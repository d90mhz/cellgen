VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

LAYER POLY1
  TYPE	MASTERSLICE ;
END POLY1

LAYER METAL1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.72  ;
  WIDTH		0.23 ;
  SPACING	0.23 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 0.00013153 ;
  EDGECAPACITANCE 8.7703e-05 ;
  CURRENTDEN 0 ;
END METAL1

LAYER VIA12
  TYPE	CUT ;
END VIA12

LAYER METAL2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.72  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 7.0018e-05 ;
  EDGECAPACITANCE 8.3115e-05 ;
  CURRENTDEN 0 ;
END METAL2

LAYER VIA23
  TYPE	CUT ;
END VIA23

LAYER METAL3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.72  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 6.3069e-05 ;
  EDGECAPACITANCE 0.00010028 ;
  CURRENTDEN 0 ;
END METAL3

LAYER VIA34
  TYPE	CUT ;
END VIA34

LAYER METAL4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.72  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 5.9911e-05 ;
  EDGECAPACITANCE 8.2087e-05 ;
  CURRENTDEN 0 ;
END METAL4

LAYER VIA45
  TYPE	CUT ;
END VIA45

LAYER METAL5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.12  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 4.8201e-05 ;
  EDGECAPACITANCE 5.7592e-05 ;
  CURRENTDEN 0 ;
END METAL5

LAYER VIA56
  TYPE	CUT ;
END VIA56

LAYER METAL6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.32  ;
  WIDTH		0.44 ;
  SPACING	0.46 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.045 ;
  CAPACITANCE	CPERSQDIST 2.5892e-05 ;
  EDGECAPACITANCE 8.5718e-05 ;
  CURRENTDEN 0 ;
END METAL6

LAYER OVERLAP
  TYPE	OVERLAP ;
END OVERLAP

LAYER NWELL
  TYPE	MASTERSLICE ;
END NWELL

LAYER DIFF
  TYPE	MASTERSLICE ;
END DIFF

LAYER PDIFF
  TYPE	MASTERSLICE ;
END PDIFF

LAYER PIMP
  TYPE	MASTERSLICE ;
END PIMP

LAYER P2V
  TYPE	MASTERSLICE ;
END P2V

LAYER NDIFF
  TYPE	MASTERSLICE ;
END NDIFF

LAYER NIMP
  TYPE	MASTERSLICE ;
END NIMP

LAYER N2V
  TYPE	MASTERSLICE ;
END N2V

LAYER CONT
  TYPE	MASTERSLICE ;
END CONT

SPACING
  SAMENET METAL1  METAL1	0.23 ;
  SAMENET METAL2  METAL2	0.28 ;
  SAMENET METAL3  METAL3	0.28 ;
  SAMENET METAL4  METAL4	0.28 ;
  SAMENET METAL5  METAL5	0.28 ;
  SAMENET METAL6  METAL6	0.46 ;
  SAMENET VIA12  VIA12	0.26 ;
  SAMENET VIA23  VIA23	0.26 ;
  SAMENET VIA34  VIA34	0.26 ;
  SAMENET VIA45  VIA45	0.26 ;
  SAMENET VIA56  VIA56	0.35 ;
END SPACING

VIA via5 DEFAULT
  LAYER METAL5 ;
    RECT -0.240 -0.190 0.240 0.190 ;
  LAYER VIA56 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER METAL6 ;
    RECT -0.270 -0.270 0.270 0.270 ;
  RESISTANCE 2.54 ;
END via5

VIA via4 DEFAULT
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL5 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via4

VIA via3_2 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.535 0.140 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via3_2

VIA via3_1 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL3 ;
    RECT -0.535 -0.140 0.190 0.140 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via3_1

VIA via3 DEFAULT
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via3

VIA via2_2 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL2 ;
    RECT -0.190 -0.140 0.190 0.395 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via2_2

VIA via2_1 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL2 ;
    RECT -0.190 -0.395 0.190 0.140 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via2_1

VIA via2 DEFAULT
  LAYER METAL2 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via2

VIA via1 DEFAULT
  LAYER METAL1 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL2 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via1


VIARULE via1Array GENERATE
  LAYER METAL1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA12 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via1Array

VIARULE via2Array GENERATE
  LAYER METAL3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA23 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via2Array

VIARULE via3Array GENERATE
  LAYER METAL3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA34 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER METAL5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA45 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER METAL5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.09 ;
    METALOVERHANG 0 ;
  LAYER VIA56 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.71 BY 0.71 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER METAL1 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER METAL2 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER METAL3 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER METAL4 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER METAL5 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER METAL6 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL6 ;
    DIRECTION VERTICAL ;
END TURNM6

SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 X Y ;
    SIZE	235.000 BY 235.000 ;
END  corner

SITE  pad
    CLASS	PAD ;
    SYMMETRY	R90 X Y ;
    SIZE	0.100 BY 235.000 ;
END  pad

SITE  tsm3site
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	7.20 BY 5.04 ;
END  tsm3site

SITE  CoreSite
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	7.20 BY 5.04 ;
END  CoreSite
