VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

LAYER POLY1
  TYPE	MASTERSLICE ;
END POLY1

LAYER METAL1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.72  ;
  WIDTH		0.23 ;
  SPACING	0.23 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 0.00013153 ;
  EDGECAPACITANCE 8.7703e-05 ;
  CURRENTDEN 0 ;
END METAL1

LAYER VIA12
  TYPE	CUT ;
END VIA12

LAYER METAL2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.72  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 7.0018e-05 ;
  EDGECAPACITANCE 8.3115e-05 ;
  CURRENTDEN 0 ;
END METAL2

LAYER VIA23
  TYPE	CUT ;
END VIA23

LAYER METAL3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.72  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 6.3069e-05 ;
  EDGECAPACITANCE 0.00010028 ;
  CURRENTDEN 0 ;
END METAL3

LAYER VIA34
  TYPE	CUT ;
END VIA34

LAYER METAL4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.72  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 5.9911e-05 ;
  EDGECAPACITANCE 8.2087e-05 ;
  CURRENTDEN 0 ;
END METAL4

LAYER VIA45
  TYPE	CUT ;
END VIA45

LAYER METAL5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.12  ;
  WIDTH		0.28 ;
  SPACING	0.28 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 4.8201e-05 ;
  EDGECAPACITANCE 5.7592e-05 ;
  CURRENTDEN 0 ;
END METAL5

LAYER VIA56
  TYPE	CUT ;
END VIA56

LAYER METAL6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.32  ;
  WIDTH		0.44 ;
  SPACING	0.46 ;
  SPACING	0.6 RANGE 10 100000 ;
  RESISTANCE	RPERSQ 0.045 ;
  CAPACITANCE	CPERSQDIST 2.5892e-05 ;
  EDGECAPACITANCE 8.5718e-05 ;
  CURRENTDEN 0 ;
END METAL6

LAYER OVERLAP
  TYPE	OVERLAP ;
END OVERLAP

LAYER NWELL
  TYPE	MASTERSLICE ;
END NWELL

LAYER DIFF
  TYPE	MASTERSLICE ;
END DIFF

LAYER PDIFF
  TYPE	MASTERSLICE ;
END PDIFF

LAYER PIMP
  TYPE	MASTERSLICE ;
END PIMP

LAYER P2V
  TYPE	MASTERSLICE ;
END P2V

LAYER NDIFF
  TYPE	MASTERSLICE ;
END NDIFF

LAYER NIMP
  TYPE	MASTERSLICE ;
END NIMP

LAYER N2V
  TYPE	MASTERSLICE ;
END N2V

LAYER CONT
  TYPE	MASTERSLICE ;
END CONT

SPACING
  SAMENET METAL1  METAL1	0.23 ;
  SAMENET METAL2  METAL2	0.28 ;
  SAMENET METAL3  METAL3	0.28 ;
  SAMENET METAL4  METAL4	0.28 ;
  SAMENET METAL5  METAL5	0.28 ;
  SAMENET METAL6  METAL6	0.46 ;
  SAMENET VIA12  VIA12	0.26 ;
  SAMENET VIA23  VIA23	0.26 ;
  SAMENET VIA34  VIA34	0.26 ;
  SAMENET VIA45  VIA45	0.26 ;
  SAMENET VIA56  VIA56	0.35 ;
END SPACING

VIA via5 DEFAULT
  LAYER METAL5 ;
    RECT -0.240 -0.190 0.240 0.190 ;
  LAYER VIA56 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER METAL6 ;
    RECT -0.270 -0.270 0.270 0.270 ;
  RESISTANCE 2.54 ;
END via5

VIA via4 DEFAULT
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL5 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via4

VIA via3_2 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.535 0.140 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via3_2

VIA via3_1 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL3 ;
    RECT -0.535 -0.140 0.190 0.140 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via3_1

VIA via3 DEFAULT
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL4 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via3

VIA via2_2 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL2 ;
    RECT -0.190 -0.140 0.190 0.395 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via2_2

VIA via2_1 DEFAULT
  TOPOFSTACKONLY
  LAYER METAL2 ;
    RECT -0.190 -0.395 0.190 0.140 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via2_1

VIA via2 DEFAULT
  LAYER METAL2 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL3 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via2

VIA via1 DEFAULT
  LAYER METAL1 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
  LAYER METAL2 ;
    RECT -0.190 -0.140 0.190 0.140 ;
  RESISTANCE 6.40 ;
END via1


VIARULE via1Array GENERATE
  LAYER METAL1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA12 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via1Array

VIARULE via2Array GENERATE
  LAYER METAL3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA23 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via2Array

VIARULE via3Array GENERATE
  LAYER METAL3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA34 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER METAL5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER VIA45 ;
    RECT -0.13 -0.13 0.13 0.13 ;
    SPACING 0.52 BY 0.52 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER METAL5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.06 ;
    METALOVERHANG 0 ;
  LAYER METAL6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.09 ;
    METALOVERHANG 0 ;
  LAYER VIA56 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.71 BY 0.71 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER METAL1 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER METAL2 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER METAL3 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER METAL4 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER METAL5 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER METAL6 ;
    DIRECTION HORIZONTAL ;
  LAYER METAL6 ;
    DIRECTION VERTICAL ;
END TURNM6

SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 X Y ;
    SIZE	235.000 BY 235.000 ;
END  corner

SITE  pad
    CLASS	PAD ;
    SYMMETRY	R90 X Y ;
    SIZE	0.100 BY 235.000 ;
END  pad

SITE  tsm3site
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	7.20 BY 5.04 ;
END  tsm3site

SITE  CoreSite
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	7.20 BY 5.04 ;
END  CoreSite
SITE  TDCoverSite
    CLASS       CORE ;
    SIZE        1.000 BY 1.000 ;
END  TDCoverSite

SITE  SBlockSite
    CLASS       CORE ;
    SIZE        1.000 BY 1.000 ;
END  SBlockSite

SITE  PortCellSite
    CLASS       PAD ;
    SIZE        1.000 BY 1.000 ;
END  PortCellSite

SITE  Core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SIZE        8.000 BY 5.040 ;
END  Core

MACRO inv_1
  CLASS CORE ;
  FOREIGN inv_1 -0.360 -2.270 ;
  ORIGIN 0.360 2.270 ;
  SIZE 4.320 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -0.360 2.370 3.960 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -0.360 -2.670 3.960 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.580 -0.060 0.865 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in0
  OBS
    LAYER NWELL ;
    RECT -1.080 0.000 4.680 3.310 ;
    LAYER NIMP ;
    RECT -0.390 -1.725 3.990 0.000 ;
    RECT -0.460 2.225 4.060 2.990 ;
    LAYER PIMP ;
    RECT -0.390 0.000 2.550 2.225 ;
    RECT -0.460 -2.490 4.060 -1.725 ;
    LAYER N2V ;
    RECT -0.390 -1.725 3.990 0.000 ;
    LAYER P2V ;
    RECT -0.390 0.000 2.550 2.225 ;
    LAYER DIFF ;
    RECT -0.360 2.325 3.960 2.880 ;
    RECT -0.210 -1.325 3.810 -0.485 ;
    RECT -0.360 -2.380 3.960 -1.825 ;
    RECT -0.210 0.450 2.370 1.850 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.070 ;
    RECT 0.990 0.000 1.170 2.070 ;
    RECT 0.270 -0.330 1.170 0.330 ;
    RECT 1.710 0.000 1.890 2.070 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT 0.270 -1.545 0.450 0.000 ;
    RECT 0.990 -1.545 1.170 0.000 ;
    RECT 0.270 -0.330 1.170 0.330 ;
    RECT 1.710 -1.545 1.890 0.000 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT 2.430 -1.545 2.610 0.000 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT 3.150 -1.545 3.330 0.000 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    LAYER METAL1 ;
    RECT -0.360 2.370 3.960 3.170 ;
    RECT -0.360 -2.670 3.960 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.535 -0.010 0.915 0.270 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.000 0.835 1.150 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT 1.325 1.150 1.555 2.770 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT 2.045 0.000 2.275 1.150 ;
    RECT 0.605 -0.090 2.275 0.140 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT -0.115 -2.270 0.115 -0.905 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 0.000 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT 1.325 -2.270 1.555 -0.905 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT 2.045 -0.905 2.275 0.000 ;
    RECT 0.605 -0.090 2.275 0.140 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT 2.765 -2.270 2.995 -0.905 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT 3.485 -0.905 3.715 0.000 ;
    RECT 2.045 -0.090 3.715 0.140 ;
    LAYER METAL2 ;
    RECT 0.580 -0.060 0.865 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    LAYER VIA12 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.595 0.000 0.855 0.260 ;
  END
END inv_1
MACRO nand2_1
  CLASS CORE ;
  FOREIGN nand2_1 -3.240 -2.270 ;
  ORIGIN 3.240 2.270 ;
  SIZE 7.920 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.240 2.370 4.680 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.240 -2.670 4.680 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 1.300 -0.060 1.585 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in1
  OBS
    LAYER NWELL ;
    RECT -3.960 0.000 5.400 3.310 ;
    LAYER NIMP ;
    RECT -3.270 -1.725 4.710 0.000 ;
    RECT -3.340 2.225 4.780 2.990 ;
    LAYER PIMP ;
    RECT -1.830 0.000 3.270 2.225 ;
    RECT -3.340 -2.490 4.780 -1.725 ;
    LAYER N2V ;
    RECT -3.270 -1.725 4.710 0.000 ;
    LAYER P2V ;
    RECT -1.830 0.000 3.270 2.225 ;
    LAYER DIFF ;
    RECT -3.240 2.325 4.680 2.880 ;
    RECT -3.090 -1.325 4.530 -0.485 ;
    RECT -3.240 -2.380 4.680 -1.825 ;
    RECT -1.650 0.450 3.090 1.850 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.070 ;
    RECT 0.990 0.000 1.170 2.070 ;
    RECT -0.450 0.000 -0.270 2.070 ;
    RECT 1.710 0.000 1.890 2.070 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.070 ;
    RECT 2.430 0.000 2.610 2.070 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT 0.270 -1.545 0.450 0.000 ;
    RECT 0.990 -1.545 1.170 0.000 ;
    RECT -0.450 -1.545 -0.270 0.000 ;
    RECT 1.710 -1.545 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.545 -0.990 0.000 ;
    RECT 2.430 -1.545 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 -1.545 -1.710 0.000 ;
    RECT 3.150 -1.545 3.330 0.000 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 -1.545 -2.430 0.000 ;
    RECT 3.870 -1.545 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    LAYER METAL1 ;
    RECT -3.240 2.370 4.680 3.170 ;
    RECT -3.240 -2.670 4.680 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 1.255 -0.010 1.635 0.270 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 1.150 0.835 2.770 ;
    RECT 0.605 1.150 0.835 2.770 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 0.565 0.115 1.150 ;
    RECT 1.325 0.000 1.555 1.150 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 1.150 -0.605 2.770 ;
    RECT 2.045 1.150 2.275 2.770 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT -1.555 0.565 -1.325 1.150 ;
    RECT 2.765 0.000 2.995 1.150 ;
    RECT -1.555 0.565 0.115 0.795 ;
    RECT 1.325 -0.010 2.995 0.220 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -1.630 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -2.270 0.115 -0.905 ;
    RECT 1.325 -0.905 1.555 0.000 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -0.905 -0.605 -0.330 ;
    RECT 2.045 -1.630 2.275 -0.905 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -1.630 2.275 -1.400 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -2.270 -1.325 -0.905 ;
    RECT 2.765 -0.905 2.995 0.000 ;
    RECT 1.325 -0.010 2.995 0.220 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -2.275 -0.905 -2.045 -0.330 ;
    RECT 3.485 -1.630 3.715 -0.905 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT 2.045 -1.630 3.715 -1.400 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -2.270 -2.765 -0.905 ;
    RECT 4.205 -0.905 4.435 0.000 ;
    RECT 2.765 -0.010 4.435 0.220 ;
    LAYER METAL2 ;
    RECT 1.300 -0.060 1.585 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    LAYER VIA12 ;
    RECT 1.315 0.000 1.575 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
  END
END nand2_1
MACRO nand3_1
  CLASS CORE ;
  FOREIGN nand3_1 -3.240 -2.270 ;
  ORIGIN 3.240 2.270 ;
  SIZE 11.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.240 2.370 8.280 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.240 -2.670 8.280 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.155 -0.010 4.535 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in2
  OBS
    LAYER NWELL ;
    RECT -3.960 0.000 9.000 3.310 ;
    LAYER NIMP ;
    RECT -3.270 -1.725 8.310 0.000 ;
    RECT -3.340 2.225 8.380 2.990 ;
    LAYER PIMP ;
    RECT -1.830 0.000 6.870 2.225 ;
    RECT -3.340 -2.490 8.380 -1.725 ;
    LAYER N2V ;
    RECT -3.270 -1.725 8.310 0.000 ;
    LAYER P2V ;
    RECT -1.830 0.000 6.870 2.225 ;
    LAYER DIFF ;
    RECT -3.240 2.325 8.280 2.880 ;
    RECT -3.090 -1.325 4.530 -0.485 ;
    RECT 4.110 -1.325 8.130 -0.485 ;
    RECT -3.240 -2.380 8.280 -1.825 ;
    RECT -1.650 0.450 6.690 1.850 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.070 ;
    RECT 0.990 0.000 1.170 2.070 ;
    RECT -0.450 0.000 -0.270 2.070 ;
    RECT 1.710 0.000 1.890 2.070 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.070 ;
    RECT 2.430 0.000 2.610 2.070 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT 0.270 -1.545 0.450 0.000 ;
    RECT 0.990 -1.545 1.170 0.000 ;
    RECT -0.450 -1.545 -0.270 0.000 ;
    RECT 1.710 -1.545 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.545 -0.990 0.000 ;
    RECT 2.430 -1.545 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 -1.545 -1.710 0.000 ;
    RECT 3.150 -1.545 3.330 0.000 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 -1.545 -2.430 0.000 ;
    RECT 3.870 -1.545 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT 4.590 0.000 4.770 2.070 ;
    RECT 5.310 0.000 5.490 2.070 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT 6.030 0.000 6.210 2.070 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT 4.590 -1.545 4.770 0.000 ;
    RECT 5.310 -1.545 5.490 0.000 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT 6.030 -1.545 6.210 0.000 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT 6.750 -1.545 6.930 0.000 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT 7.470 -1.545 7.650 0.000 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT 4.300 -0.130 4.720 0.290 ;
    LAYER METAL1 ;
    RECT -3.240 2.370 8.280 3.170 ;
    RECT -3.240 -2.670 8.280 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 4.155 -0.100 4.625 0.335 ;
    RECT 4.855 -0.010 5.235 0.270 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT 2.765 0.565 4.435 0.795 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 1.150 0.835 2.770 ;
    RECT 0.605 1.150 0.835 2.770 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 0.565 0.115 1.150 ;
    RECT 1.325 0.565 1.555 1.150 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 1.150 -0.605 2.770 ;
    RECT 2.045 1.150 2.275 2.770 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT -1.555 0.565 -1.325 1.150 ;
    RECT 2.765 0.565 2.995 1.150 ;
    RECT -1.555 0.565 0.115 0.795 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT 4.205 0.565 4.435 1.150 ;
    RECT 2.765 0.565 5.155 0.795 ;
    RECT 4.925 0.000 5.155 0.795 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT 4.925 1.150 5.155 2.770 ;
    RECT 5.590 1.035 5.930 1.265 ;
    RECT 4.925 -0.010 5.875 0.220 ;
    RECT 5.645 0.000 5.875 1.150 ;
    RECT 6.310 1.035 6.650 1.265 ;
    RECT 6.365 1.150 6.595 2.770 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -1.630 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.325 -0.905 1.555 -0.330 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -2.270 0.115 -0.905 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -0.905 -0.605 -0.330 ;
    RECT 2.045 -1.630 2.275 -0.905 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -1.630 2.275 -1.400 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.765 -0.905 2.995 -0.330 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT -1.555 -2.270 -1.325 -0.905 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -2.275 -0.905 -2.045 -0.330 ;
    RECT 3.485 -1.630 3.715 -0.905 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT 2.045 -1.630 3.715 -1.400 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT -2.995 -2.270 -2.765 -0.905 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT 4.205 -1.630 4.435 -0.905 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT 4.925 -0.905 5.155 0.000 ;
    RECT 5.590 -1.020 5.930 -0.790 ;
    RECT 5.645 -1.630 5.875 -0.905 ;
    RECT 4.205 -1.630 5.875 -1.400 ;
    RECT 6.310 -1.020 6.650 -0.790 ;
    RECT 6.365 -0.905 6.595 0.000 ;
    RECT 4.925 -0.010 6.595 0.220 ;
    RECT 7.030 -1.020 7.370 -0.790 ;
    RECT 7.085 -1.630 7.315 -0.905 ;
    RECT 5.645 -1.630 7.315 -1.400 ;
    RECT 7.750 -1.020 8.090 -0.790 ;
    RECT 7.805 -0.905 8.035 0.000 ;
    RECT 6.365 -0.010 8.035 0.220 ;
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT 4.155 -0.010 4.535 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 4.400 -0.030 4.620 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT 5.650 2.425 5.870 2.645 ;
    RECT 5.650 -2.145 5.870 -1.925 ;
    RECT 6.370 2.425 6.590 2.645 ;
    RECT 6.370 -2.145 6.590 -1.925 ;
    RECT 7.090 2.425 7.310 2.645 ;
    RECT 7.090 -2.145 7.310 -1.925 ;
    RECT 7.810 2.425 8.030 2.645 ;
    RECT 7.810 -2.145 8.030 -1.925 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    RECT 5.650 1.040 5.870 1.260 ;
    RECT 6.370 1.040 6.590 1.260 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT 4.930 -1.015 5.150 -0.795 ;
    RECT 5.650 -1.015 5.870 -0.795 ;
    RECT 6.370 -1.015 6.590 -0.795 ;
    RECT 7.090 -1.015 7.310 -0.795 ;
    RECT 7.810 -1.015 8.030 -0.795 ;
    LAYER VIA12 ;
    RECT 4.915 0.000 5.175 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT 4.215 0.000 4.475 0.260 ;
  END
END nand3_1
MACRO nand4_1
  CLASS CORE ;
  FOREIGN nand4_1 -6.840 -2.270 ;
  ORIGIN 6.840 2.270 ;
  SIZE 15.120 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -6.840 2.370 8.280 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -6.840 -2.670 8.280 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.155 -0.010 4.535 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in2
  PIN in3
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -3.765 -0.010 -3.385 0.270 ;
    END
  END in3
  OBS
    LAYER NWELL ;
    RECT -7.560 0.000 9.000 3.310 ;
    LAYER NIMP ;
    RECT -6.870 -1.725 8.310 0.000 ;
    RECT -6.940 2.225 8.380 2.990 ;
    LAYER PIMP ;
    RECT -5.430 0.000 6.870 2.225 ;
    RECT -6.940 -2.490 8.380 -1.725 ;
    LAYER N2V ;
    RECT -6.870 -1.725 8.310 0.000 ;
    LAYER P2V ;
    RECT -5.430 0.000 6.870 2.225 ;
    LAYER DIFF ;
    RECT -6.840 2.325 8.280 2.880 ;
    RECT -3.090 -1.325 4.530 -0.485 ;
    RECT 4.110 -1.325 8.130 -0.485 ;
    RECT -6.690 -1.325 -2.670 -0.485 ;
    RECT -6.840 -2.380 8.280 -1.825 ;
    RECT -5.250 0.450 6.690 1.850 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.070 ;
    RECT 0.990 0.000 1.170 2.070 ;
    RECT -0.450 0.000 -0.270 2.070 ;
    RECT 1.710 0.000 1.890 2.070 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.070 ;
    RECT 2.430 0.000 2.610 2.070 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT 0.270 -1.545 0.450 0.000 ;
    RECT 0.990 -1.545 1.170 0.000 ;
    RECT -0.450 -1.545 -0.270 0.000 ;
    RECT 1.710 -1.545 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.545 -0.990 0.000 ;
    RECT 2.430 -1.545 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 -1.545 -1.710 0.000 ;
    RECT 3.150 -1.545 3.330 0.000 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 -1.545 -2.430 0.000 ;
    RECT 3.870 -1.545 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 0.000 -3.150 2.070 ;
    RECT 4.590 0.000 4.770 2.070 ;
    RECT -4.050 0.000 -3.870 2.070 ;
    RECT 5.310 0.000 5.490 2.070 ;
    RECT -4.050 -0.330 -3.150 0.330 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT -4.770 0.000 -4.590 2.070 ;
    RECT 6.030 0.000 6.210 2.070 ;
    RECT -4.770 -0.330 -3.870 0.330 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT -3.330 -1.545 -3.150 0.000 ;
    RECT 4.590 -1.545 4.770 0.000 ;
    RECT -4.050 -1.545 -3.870 0.000 ;
    RECT 5.310 -1.545 5.490 0.000 ;
    RECT -4.050 -0.330 -3.150 0.330 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT -4.770 -1.545 -4.590 0.000 ;
    RECT 6.030 -1.545 6.210 0.000 ;
    RECT -4.770 -0.330 -3.870 0.330 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT -5.490 -1.545 -5.310 0.000 ;
    RECT 6.750 -1.545 6.930 0.000 ;
    RECT -5.490 -0.330 -4.590 0.330 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT -6.210 -1.545 -6.030 0.000 ;
    RECT 7.470 -1.545 7.650 0.000 ;
    RECT -6.210 -0.330 -5.310 0.330 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT 4.300 -0.130 4.720 0.290 ;
    RECT -3.620 -0.130 -3.200 0.290 ;
    LAYER METAL1 ;
    RECT -6.840 2.370 8.280 3.170 ;
    RECT -6.840 -2.670 8.280 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 4.155 -0.100 4.625 0.335 ;
    RECT -3.765 -0.100 -3.295 0.335 ;
    RECT 4.855 -0.010 5.235 0.270 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -1.555 0.565 0.115 0.795 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT -2.995 0.565 -1.325 0.795 ;
    RECT 2.765 0.565 4.435 0.795 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 1.150 0.835 2.770 ;
    RECT 0.605 1.150 0.835 2.770 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 0.565 0.115 1.150 ;
    RECT 1.325 0.565 1.555 1.150 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -0.115 0.565 1.555 0.795 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 1.150 -0.605 2.770 ;
    RECT 2.045 1.150 2.275 2.770 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT -1.555 0.565 -1.325 1.150 ;
    RECT 2.765 0.565 2.995 1.150 ;
    RECT -1.555 0.565 0.115 0.795 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT -3.050 1.035 -2.710 1.265 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT -2.995 0.565 -2.765 1.150 ;
    RECT 4.205 0.565 4.435 1.150 ;
    RECT -2.995 0.565 -1.325 0.795 ;
    RECT 2.765 0.565 5.155 0.795 ;
    RECT 4.925 0.000 5.155 0.795 ;
    RECT -3.770 1.035 -3.430 1.265 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT -3.715 1.150 -3.485 2.770 ;
    RECT 4.925 1.150 5.155 2.770 ;
    RECT -4.490 1.035 -4.150 1.265 ;
    RECT 5.590 1.035 5.930 1.265 ;
    RECT -4.435 0.565 -2.765 0.795 ;
    RECT 4.925 -0.010 5.875 0.220 ;
    RECT -4.435 0.565 -4.205 1.150 ;
    RECT 5.645 0.000 5.875 1.150 ;
    RECT -5.210 1.035 -4.870 1.265 ;
    RECT 6.310 1.035 6.650 1.265 ;
    RECT -5.155 1.150 -4.925 2.770 ;
    RECT 6.365 1.150 6.595 2.770 ;
    RECT -1.555 -1.630 0.115 -1.400 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT -2.995 -1.630 -1.325 -1.400 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -1.630 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -1.630 0.115 -0.905 ;
    RECT 1.325 -0.905 1.555 -0.330 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -0.905 -0.605 -0.330 ;
    RECT 2.045 -1.630 2.275 -0.905 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -1.630 2.275 -1.400 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -1.630 -1.325 -0.905 ;
    RECT 2.765 -0.905 2.995 -0.330 ;
    RECT -1.555 -1.630 0.115 -1.400 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -2.275 -0.905 -2.045 -0.330 ;
    RECT 3.485 -1.630 3.715 -0.905 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT 2.045 -1.630 3.715 -1.400 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -1.630 -2.765 -0.905 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT -2.995 -1.630 -1.325 -1.400 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -0.905 -2.765 -0.330 ;
    RECT 4.205 -1.630 4.435 -0.905 ;
    RECT -2.995 -1.630 -1.325 -1.400 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT -2.995 -1.630 -2.765 -0.905 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT -3.770 -1.020 -3.430 -0.790 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT -3.715 -2.270 -3.485 -0.905 ;
    RECT 4.925 -0.905 5.155 0.000 ;
    RECT -4.490 -1.020 -4.150 -0.790 ;
    RECT 5.590 -1.020 5.930 -0.790 ;
    RECT -4.435 -0.905 -4.205 -0.330 ;
    RECT 5.645 -1.630 5.875 -0.905 ;
    RECT -4.435 -0.560 -2.765 -0.330 ;
    RECT 4.205 -1.630 5.875 -1.400 ;
    RECT -5.210 -1.020 -4.870 -0.790 ;
    RECT 6.310 -1.020 6.650 -0.790 ;
    RECT -5.155 -2.270 -4.925 -0.905 ;
    RECT 6.365 -0.905 6.595 0.000 ;
    RECT 4.925 -0.010 6.595 0.220 ;
    RECT -5.930 -1.020 -5.590 -0.790 ;
    RECT 7.030 -1.020 7.370 -0.790 ;
    RECT -5.875 -0.905 -5.645 -0.330 ;
    RECT 7.085 -1.630 7.315 -0.905 ;
    RECT -5.875 -0.560 -4.205 -0.330 ;
    RECT 5.645 -1.630 7.315 -1.400 ;
    RECT -6.650 -1.020 -6.310 -0.790 ;
    RECT 7.750 -1.020 8.090 -0.790 ;
    RECT -6.595 -2.270 -6.365 -0.905 ;
    RECT 7.805 -0.905 8.035 0.000 ;
    RECT 6.365 -0.010 8.035 0.220 ;
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT 4.155 -0.010 4.535 0.270 ;
    RECT -3.765 -0.010 -3.385 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 4.400 -0.030 4.620 0.190 ;
    RECT -3.520 -0.030 -3.300 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT -3.710 2.425 -3.490 2.645 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT -3.710 -2.145 -3.490 -1.925 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT -4.430 2.425 -4.210 2.645 ;
    RECT 5.650 2.425 5.870 2.645 ;
    RECT -4.430 -2.145 -4.210 -1.925 ;
    RECT 5.650 -2.145 5.870 -1.925 ;
    RECT -5.150 2.425 -4.930 2.645 ;
    RECT 6.370 2.425 6.590 2.645 ;
    RECT -5.150 -2.145 -4.930 -1.925 ;
    RECT 6.370 -2.145 6.590 -1.925 ;
    RECT -5.870 2.425 -5.650 2.645 ;
    RECT 7.090 2.425 7.310 2.645 ;
    RECT -5.870 -2.145 -5.650 -1.925 ;
    RECT 7.090 -2.145 7.310 -1.925 ;
    RECT -6.590 2.425 -6.370 2.645 ;
    RECT 7.810 2.425 8.030 2.645 ;
    RECT -6.590 -2.145 -6.370 -1.925 ;
    RECT 7.810 -2.145 8.030 -1.925 ;
    RECT -2.990 1.040 -2.770 1.260 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT -3.710 1.040 -3.490 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    RECT -4.430 1.040 -4.210 1.260 ;
    RECT 5.650 1.040 5.870 1.260 ;
    RECT -5.150 1.040 -4.930 1.260 ;
    RECT 6.370 1.040 6.590 1.260 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT -3.710 -1.015 -3.490 -0.795 ;
    RECT 4.930 -1.015 5.150 -0.795 ;
    RECT -4.430 -1.015 -4.210 -0.795 ;
    RECT 5.650 -1.015 5.870 -0.795 ;
    RECT -5.150 -1.015 -4.930 -0.795 ;
    RECT 6.370 -1.015 6.590 -0.795 ;
    RECT -5.870 -1.015 -5.650 -0.795 ;
    RECT 7.090 -1.015 7.310 -0.795 ;
    RECT -6.590 -1.015 -6.370 -0.795 ;
    RECT 7.810 -1.015 8.030 -0.795 ;
    LAYER VIA12 ;
    RECT 4.915 0.000 5.175 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT 4.215 0.000 4.475 0.260 ;
    RECT -3.705 0.000 -3.445 0.260 ;
  END
END nand4_1
MACRO nor2_1
  CLASS CORE ;
  FOREIGN nor2_1 -0.360 -2.270 ;
  ORIGIN 0.360 2.270 ;
  SIZE 2.160 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -0.360 2.370 1.800 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -0.360 -2.670 1.800 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 1.300 -0.060 1.585 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in1
  OBS
    LAYER NWELL ;
    RECT -1.080 0.000 2.520 3.310 ;
    LAYER NIMP ;
    RECT -0.390 -1.725 1.830 0.000 ;
    RECT -0.460 2.225 1.900 2.990 ;
    LAYER PIMP ;
    RECT -0.390 0.000 1.830 2.225 ;
    RECT -0.460 -2.490 1.900 -1.725 ;
    LAYER N2V ;
    RECT -0.390 -1.725 1.830 0.000 ;
    LAYER P2V ;
    RECT -0.390 0.000 1.830 2.225 ;
    LAYER DIFF ;
    RECT -0.360 2.325 1.800 2.880 ;
    RECT -0.210 -1.115 1.650 -0.695 ;
    RECT -0.360 -2.380 1.800 -1.825 ;
    RECT -0.210 0.940 1.650 1.360 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 1.580 ;
    RECT 0.990 0.000 1.170 1.580 ;
    RECT 0.270 -1.335 0.450 0.000 ;
    RECT 0.990 -1.335 1.170 0.000 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    LAYER METAL1 ;
    RECT -0.360 2.370 1.800 3.170 ;
    RECT -0.360 -2.670 1.800 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 1.255 -0.010 1.635 0.270 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -2.270 0.835 -0.905 ;
    RECT 0.605 -2.270 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -0.905 0.115 -0.330 ;
    RECT 1.325 -0.905 1.555 0.000 ;
    RECT -0.115 -0.560 1.555 -0.330 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT 1.325 0.000 1.555 1.150 ;
    LAYER METAL2 ;
    RECT 1.300 -0.060 1.585 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    LAYER VIA12 ;
    RECT 1.315 0.000 1.575 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
  END
END nor2_1
MACRO nor3_1
  CLASS CORE ;
  FOREIGN nor3_1 -3.240 -2.270 ;
  ORIGIN 3.240 2.270 ;
  SIZE 11.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.240 2.370 8.280 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.240 -2.670 8.280 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.155 -0.010 4.535 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in2
  OBS
    LAYER NWELL ;
    RECT -3.960 0.000 9.000 3.310 ;
    LAYER NIMP ;
    RECT -3.270 -1.725 8.310 0.000 ;
    RECT -3.340 2.225 8.380 2.990 ;
    LAYER PIMP ;
    RECT -1.830 0.000 6.870 2.225 ;
    RECT -3.340 -2.490 8.380 -1.725 ;
    LAYER N2V ;
    RECT -3.270 -1.725 8.310 0.000 ;
    LAYER P2V ;
    RECT -1.830 0.000 6.870 2.225 ;
    LAYER DIFF ;
    RECT -3.240 2.325 8.280 2.880 ;
    RECT -3.090 -1.325 8.130 -0.485 ;
    RECT -3.240 -2.380 8.280 -1.825 ;
    RECT 4.110 0.450 6.690 1.850 ;
    RECT -1.650 0.450 4.530 1.850 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.070 ;
    RECT 0.990 0.000 1.170 2.070 ;
    RECT -0.450 0.000 -0.270 2.070 ;
    RECT 1.710 0.000 1.890 2.070 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.070 ;
    RECT 2.430 0.000 2.610 2.070 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT 0.270 -1.545 0.450 0.000 ;
    RECT 0.990 -1.545 1.170 0.000 ;
    RECT -0.450 -1.545 -0.270 0.000 ;
    RECT 1.710 -1.545 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.545 -0.990 0.000 ;
    RECT 2.430 -1.545 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 -1.545 -1.710 0.000 ;
    RECT 3.150 -1.545 3.330 0.000 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 -1.545 -2.430 0.000 ;
    RECT 3.870 -1.545 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT 4.590 0.000 4.770 2.070 ;
    RECT 5.310 0.000 5.490 2.070 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT 6.030 0.000 6.210 2.070 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT 4.590 -1.545 4.770 0.000 ;
    RECT 5.310 -1.545 5.490 0.000 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT 6.030 -1.545 6.210 0.000 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT 6.750 -1.545 6.930 0.000 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT 7.470 -1.545 7.650 0.000 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT 4.300 -0.130 4.720 0.290 ;
    LAYER METAL1 ;
    RECT -3.240 2.370 8.280 3.170 ;
    RECT -3.240 -2.670 8.280 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 4.155 -0.100 4.625 0.335 ;
    RECT 4.855 -0.010 5.235 0.270 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT 2.765 0.565 4.435 0.795 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT 0.605 1.150 0.835 2.130 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT 1.325 0.565 1.555 1.150 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 0.565 -0.605 1.150 ;
    RECT 2.045 1.150 2.275 2.130 ;
    RECT -0.835 0.565 0.835 0.795 ;
    RECT 0.605 1.900 2.275 2.130 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT 2.765 0.565 2.995 1.150 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT -1.555 1.150 -1.325 2.770 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT 4.205 1.150 4.435 2.130 ;
    RECT 2.765 0.565 4.435 0.795 ;
    RECT 4.205 0.565 4.435 1.150 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT 4.925 0.000 5.155 1.150 ;
    RECT 5.590 1.035 5.930 1.265 ;
    RECT 5.645 1.150 5.875 2.130 ;
    RECT 4.205 1.900 5.875 2.130 ;
    RECT 6.310 1.035 6.650 1.265 ;
    RECT 6.365 0.000 6.595 1.150 ;
    RECT 4.925 -0.010 6.595 0.220 ;
    RECT -0.115 -0.560 1.555 -0.330 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -2.270 0.835 -0.905 ;
    RECT 0.605 -2.270 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -0.905 0.115 -0.330 ;
    RECT 1.325 -0.905 1.555 -0.330 ;
    RECT -0.115 -0.560 1.555 -0.330 ;
    RECT -0.115 -0.560 1.555 -0.330 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -2.270 -0.605 -0.905 ;
    RECT 2.045 -2.270 2.275 -0.905 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -0.905 -1.325 -0.330 ;
    RECT 2.765 -0.905 2.995 -0.330 ;
    RECT -1.555 -0.560 0.115 -0.330 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -2.275 -2.270 -2.045 -0.905 ;
    RECT 3.485 -2.270 3.715 -0.905 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -0.905 -2.765 -0.330 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT -2.995 -0.560 -1.325 -0.330 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT 2.765 -0.560 5.155 -0.330 ;
    RECT 4.925 -0.560 5.155 0.000 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT 4.925 -2.270 5.155 -0.905 ;
    RECT 5.590 -1.020 5.930 -0.790 ;
    RECT 4.925 -0.010 5.875 0.220 ;
    RECT 5.645 -0.905 5.875 0.000 ;
    RECT 6.310 -1.020 6.650 -0.790 ;
    RECT 6.365 -2.270 6.595 -0.905 ;
    RECT 7.030 -1.020 7.370 -0.790 ;
    RECT 5.645 -0.010 7.315 0.220 ;
    RECT 7.085 -0.905 7.315 0.000 ;
    RECT 7.750 -1.020 8.090 -0.790 ;
    RECT 7.805 -2.270 8.035 -0.905 ;
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT 4.155 -0.010 4.535 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 4.400 -0.030 4.620 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT 5.650 2.425 5.870 2.645 ;
    RECT 5.650 -2.145 5.870 -1.925 ;
    RECT 6.370 2.425 6.590 2.645 ;
    RECT 6.370 -2.145 6.590 -1.925 ;
    RECT 7.090 2.425 7.310 2.645 ;
    RECT 7.090 -2.145 7.310 -1.925 ;
    RECT 7.810 2.425 8.030 2.645 ;
    RECT 7.810 -2.145 8.030 -1.925 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    RECT 5.650 1.040 5.870 1.260 ;
    RECT 6.370 1.040 6.590 1.260 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT 4.930 -1.015 5.150 -0.795 ;
    RECT 5.650 -1.015 5.870 -0.795 ;
    RECT 6.370 -1.015 6.590 -0.795 ;
    RECT 7.090 -1.015 7.310 -0.795 ;
    RECT 7.810 -1.015 8.030 -0.795 ;
    LAYER VIA12 ;
    RECT 4.915 0.000 5.175 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT 4.215 0.000 4.475 0.260 ;
  END
END nor3_1
MACRO aoi21_1
  CLASS CORE ;
  FOREIGN aoi21_1 -1.080 -2.270 ;
  ORIGIN 1.080 2.270 ;
  SIZE 2.880 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -1.080 2.370 1.800 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -1.080 -2.670 1.800 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 1.300 -0.060 1.585 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.885 -0.010 -0.505 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in2
  OBS
    LAYER NWELL ;
    RECT -1.800 0.000 2.520 3.310 ;
    LAYER NIMP ;
    RECT -1.110 -1.725 1.830 0.000 ;
    RECT -1.180 2.225 1.900 2.990 ;
    LAYER PIMP ;
    RECT -1.110 0.000 1.830 2.225 ;
    RECT -1.180 -2.490 1.900 -1.725 ;
    LAYER N2V ;
    RECT -1.110 -1.725 1.830 0.000 ;
    LAYER P2V ;
    RECT -1.110 0.000 1.830 2.225 ;
    LAYER DIFF ;
    RECT -1.080 -2.380 1.800 -1.825 ;
    RECT -0.210 -1.115 1.650 -0.695 ;
    RECT -0.930 -1.115 0.210 -0.695 ;
    RECT -1.080 2.325 1.800 2.880 ;
    RECT -0.930 0.940 1.650 1.360 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 1.580 ;
    RECT 0.990 0.000 1.170 1.580 ;
    RECT 0.270 -1.335 0.450 0.000 ;
    RECT 0.990 -1.335 1.170 0.000 ;
    RECT -0.450 0.000 -0.270 1.580 ;
    RECT -0.450 -1.335 -0.270 0.000 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT -0.740 -0.130 -0.320 0.290 ;
    LAYER METAL1 ;
    RECT -1.080 2.370 1.800 3.170 ;
    RECT -1.080 -2.670 1.800 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT -0.885 -0.100 -0.415 0.335 ;
    RECT 1.255 -0.010 1.635 0.270 ;
    RECT 1.325 -0.560 1.555 0.000 ;
    RECT 0.605 -0.560 1.555 -0.330 ;
    RECT 1.325 -0.115 1.555 0.115 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT 1.325 -2.270 1.555 -0.905 ;
    RECT -0.835 -2.270 -0.605 -0.905 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT 1.325 0.000 1.555 1.150 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT -0.835 0.565 -0.605 1.150 ;
    RECT -0.835 0.565 0.835 0.795 ;
    LAYER METAL2 ;
    RECT 1.300 -0.060 1.585 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT -0.885 -0.010 -0.505 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT -0.640 -0.030 -0.420 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    LAYER VIA12 ;
    RECT 1.315 0.000 1.575 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT -0.825 0.000 -0.565 0.260 ;
  END
END aoi21_1
MACRO aoi22_1
  CLASS CORE ;
  FOREIGN aoi22_1 -3.960 -2.270 ;
  ORIGIN 3.960 2.270 ;
  SIZE 9.360 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.960 2.370 5.400 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -3.960 -2.670 5.400 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -2.325 -0.010 -1.945 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in2
  PIN in3
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 2.715 -0.010 3.095 0.270 ;
    END
  END in3
  OBS
    LAYER NWELL ;
    RECT -4.680 0.000 6.120 3.310 ;
    LAYER NIMP ;
    RECT -3.990 -1.725 5.430 0.000 ;
    RECT -4.060 2.225 5.500 2.990 ;
    LAYER PIMP ;
    RECT -3.990 0.000 5.430 2.225 ;
    RECT -4.060 -2.490 5.500 -1.725 ;
    LAYER N2V ;
    RECT -3.990 -1.725 5.430 0.000 ;
    LAYER P2V ;
    RECT -3.990 0.000 5.430 2.225 ;
    LAYER DIFF ;
    RECT -3.960 -2.380 5.400 -1.825 ;
    RECT -1.650 -1.375 3.090 -0.430 ;
    RECT 2.670 -1.375 5.250 -0.430 ;
    RECT -3.810 -1.375 -1.230 -0.430 ;
    RECT -3.960 2.325 5.400 2.880 ;
    RECT -3.810 0.430 5.250 1.875 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.095 ;
    RECT 0.990 0.000 1.170 2.095 ;
    RECT -0.450 0.000 -0.270 2.095 ;
    RECT 1.710 0.000 1.890 2.095 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.095 ;
    RECT 2.430 0.000 2.610 2.095 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT 0.270 -1.595 0.450 0.000 ;
    RECT 0.990 -1.595 1.170 0.000 ;
    RECT -0.450 -1.595 -0.270 0.000 ;
    RECT 1.710 -1.595 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.595 -0.990 0.000 ;
    RECT 2.430 -1.595 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 0.000 -1.710 2.095 ;
    RECT 3.150 0.000 3.330 2.095 ;
    RECT -2.610 0.000 -2.430 2.095 ;
    RECT 3.870 0.000 4.050 2.095 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 0.000 -3.150 2.095 ;
    RECT 4.590 0.000 4.770 2.095 ;
    RECT -3.330 -0.330 -2.430 0.330 ;
    RECT 3.870 -0.330 4.770 0.330 ;
    RECT -1.890 -1.595 -1.710 0.000 ;
    RECT 3.150 -1.595 3.330 0.000 ;
    RECT -2.610 -1.595 -2.430 0.000 ;
    RECT 3.870 -1.595 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 -1.595 -3.150 0.000 ;
    RECT 4.590 -1.595 4.770 0.000 ;
    RECT -3.330 -0.330 -2.430 0.330 ;
    RECT 3.870 -0.330 4.770 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT 2.860 -0.130 3.280 0.290 ;
    RECT -2.180 -0.130 -1.760 0.290 ;
    LAYER METAL1 ;
    RECT -3.960 2.370 5.400 3.170 ;
    RECT -3.960 -2.670 5.400 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 2.715 -0.100 3.185 0.335 ;
    RECT -2.325 -0.100 -1.855 0.335 ;
    RECT 4.855 -0.010 5.235 0.270 ;
    RECT 4.925 0.000 5.155 0.795 ;
    RECT 1.325 0.565 5.155 0.795 ;
    RECT 2.045 -0.560 2.275 0.795 ;
    RECT -0.115 -1.630 1.555 -1.400 ;
    RECT -0.115 -1.630 1.555 -1.400 ;
    RECT -1.555 -1.630 0.115 -1.400 ;
    RECT 1.325 -1.630 2.995 -1.400 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -0.560 2.275 -0.330 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -1.630 0.115 -0.905 ;
    RECT 1.325 -1.630 1.555 -0.905 ;
    RECT -0.115 -1.630 1.555 -1.400 ;
    RECT -0.115 -1.630 1.555 -1.400 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -0.905 -0.605 -0.330 ;
    RECT 2.045 -0.905 2.275 -0.330 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -0.560 2.275 -0.330 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -1.630 -1.325 -0.905 ;
    RECT 2.765 -1.630 2.995 -0.905 ;
    RECT -1.555 -1.630 0.115 -1.400 ;
    RECT 1.325 -1.630 2.995 -1.400 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -0.905 -1.325 -0.330 ;
    RECT 2.765 -0.905 2.995 -0.330 ;
    RECT -1.555 -1.630 -1.325 -0.905 ;
    RECT 2.765 -1.630 2.995 -0.905 ;
    RECT -1.555 -1.630 0.115 -1.400 ;
    RECT 1.325 -1.630 2.995 -1.400 ;
    RECT -2.275 -2.270 -2.045 -0.905 ;
    RECT 3.485 -2.270 3.715 -0.905 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -0.905 -2.765 -0.330 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT -2.995 -0.560 -1.325 -0.330 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT -3.715 -2.270 -3.485 -0.905 ;
    RECT 4.925 -2.270 5.155 -0.905 ;
    RECT -3.770 -1.020 -3.430 -0.790 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT -0.835 0.565 0.835 0.795 ;
    RECT 0.605 1.900 2.275 2.130 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT 0.605 2.130 0.835 1.150 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT 1.325 0.565 1.555 1.150 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 0.565 -0.605 1.150 ;
    RECT 2.045 2.130 2.275 1.150 ;
    RECT -0.835 0.565 0.835 0.795 ;
    RECT 0.605 1.900 2.275 2.130 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT -1.555 1.150 -1.325 2.770 ;
    RECT 2.765 0.565 2.995 1.150 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT -1.555 1.150 -1.325 2.770 ;
    RECT 2.765 0.565 2.995 1.150 ;
    RECT 1.325 0.565 2.995 0.795 ;
    RECT -2.330 1.035 -1.990 1.265 ;
    RECT 3.430 1.035 3.770 1.265 ;
    RECT -2.275 0.565 -2.045 1.150 ;
    RECT 3.485 1.150 3.715 2.130 ;
    RECT -2.275 0.565 -0.605 0.795 ;
    RECT 2.045 1.900 3.715 2.130 ;
    RECT -3.050 1.035 -2.710 1.265 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT -2.995 1.150 -2.765 2.770 ;
    RECT 4.205 0.565 4.435 1.150 ;
    RECT 2.765 0.565 4.435 0.795 ;
    RECT -3.770 1.035 -3.430 1.265 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT -3.715 0.565 -3.485 1.150 ;
    RECT 4.925 1.150 5.155 2.130 ;
    RECT -3.715 0.565 -2.045 0.795 ;
    RECT 3.485 1.900 5.155 2.130 ;
    LAYER METAL2 ;
    RECT 4.900 -0.060 5.185 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT 2.715 -0.010 3.095 0.270 ;
    RECT -2.325 -0.010 -1.945 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 2.960 -0.030 3.180 0.190 ;
    RECT -2.080 -0.030 -1.860 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT -3.710 2.425 -3.490 2.645 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT -3.710 -2.145 -3.490 -1.925 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT -3.710 -1.015 -3.490 -0.795 ;
    RECT 4.930 -1.015 5.150 -0.795 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT -2.270 1.040 -2.050 1.260 ;
    RECT 3.490 1.040 3.710 1.260 ;
    RECT -2.990 1.040 -2.770 1.260 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT -3.710 1.040 -3.490 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    LAYER VIA12 ;
    RECT 4.915 0.000 5.175 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT 2.775 0.000 3.035 0.260 ;
    RECT -2.265 0.000 -2.005 0.260 ;
  END
END aoi22_1
MACRO oai21_1
  CLASS CORE ;
  FOREIGN oai21_1 -14.760 -2.270 ;
  ORIGIN 14.760 2.270 ;
  SIZE 23.040 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -14.760 2.370 8.280 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -14.760 -2.670 8.280 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 7.780 -0.060 8.065 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -8.085 -0.010 -7.705 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in2
  OBS
    LAYER NWELL ;
    RECT -15.480 0.000 9.000 3.310 ;
    LAYER NIMP ;
    RECT -14.790 -1.725 8.310 0.000 ;
    RECT -14.860 2.225 8.380 2.990 ;
    LAYER PIMP ;
    RECT -14.790 0.000 8.310 2.225 ;
    RECT -14.860 -2.490 8.380 -1.725 ;
    LAYER N2V ;
    RECT -14.790 -1.725 8.310 0.000 ;
    LAYER P2V ;
    RECT -14.790 0.000 8.310 2.225 ;
    LAYER DIFF ;
    RECT -14.760 -2.380 8.280 -1.825 ;
    RECT -6.690 0.430 8.130 1.875 ;
    RECT -14.610 0.430 -6.990 1.875 ;
    RECT -14.760 2.325 8.280 2.880 ;
    RECT -14.610 -1.375 8.130 -0.430 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.095 ;
    RECT 0.990 0.000 1.170 2.095 ;
    RECT -0.450 0.000 -0.270 2.095 ;
    RECT 1.710 0.000 1.890 2.095 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.095 ;
    RECT 2.430 0.000 2.610 2.095 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 0.000 -1.710 2.095 ;
    RECT 3.150 0.000 3.330 2.095 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 0.000 -2.430 2.095 ;
    RECT 3.870 0.000 4.050 2.095 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 0.000 -3.150 2.095 ;
    RECT 4.590 0.000 4.770 2.095 ;
    RECT -3.330 -0.330 -2.430 0.330 ;
    RECT 3.870 -0.330 4.770 0.330 ;
    RECT -4.050 0.000 -3.870 2.095 ;
    RECT 5.310 0.000 5.490 2.095 ;
    RECT -4.050 -0.330 -3.150 0.330 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT -4.770 0.000 -4.590 2.095 ;
    RECT 6.030 0.000 6.210 2.095 ;
    RECT -4.770 -0.330 -3.870 0.330 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT -5.490 0.000 -5.310 2.095 ;
    RECT 6.750 0.000 6.930 2.095 ;
    RECT -5.490 -0.330 -4.590 0.330 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT -6.210 0.000 -6.030 2.095 ;
    RECT 7.470 0.000 7.650 2.095 ;
    RECT -6.210 -0.330 -5.310 0.330 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT 0.270 -1.595 0.450 0.000 ;
    RECT 0.990 -1.595 1.170 0.000 ;
    RECT -0.450 -1.595 -0.270 0.000 ;
    RECT 1.710 -1.595 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.595 -0.990 0.000 ;
    RECT 2.430 -1.595 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 -1.595 -1.710 0.000 ;
    RECT 3.150 -1.595 3.330 0.000 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 -1.595 -2.430 0.000 ;
    RECT 3.870 -1.595 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 -1.595 -3.150 0.000 ;
    RECT 4.590 -1.595 4.770 0.000 ;
    RECT -3.330 -0.330 -2.430 0.330 ;
    RECT 3.870 -0.330 4.770 0.330 ;
    RECT -4.050 -1.595 -3.870 0.000 ;
    RECT 5.310 -1.595 5.490 0.000 ;
    RECT -4.050 -0.330 -3.150 0.330 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT -4.770 -1.595 -4.590 0.000 ;
    RECT 6.030 -1.595 6.210 0.000 ;
    RECT -4.770 -0.330 -3.870 0.330 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT -5.490 -1.595 -5.310 0.000 ;
    RECT 6.750 -1.595 6.930 0.000 ;
    RECT -5.490 -0.330 -4.590 0.330 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT -6.210 -1.595 -6.030 0.000 ;
    RECT 7.470 -1.595 7.650 0.000 ;
    RECT -6.210 -0.330 -5.310 0.330 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT -7.650 0.000 -7.470 2.095 ;
    RECT -8.370 0.000 -8.190 2.095 ;
    RECT -8.370 -0.330 -7.470 0.330 ;
    RECT -9.090 0.000 -8.910 2.095 ;
    RECT -9.090 -0.330 -8.190 0.330 ;
    RECT -9.810 0.000 -9.630 2.095 ;
    RECT -9.810 -0.330 -8.910 0.330 ;
    RECT -10.530 0.000 -10.350 2.095 ;
    RECT -10.530 -0.330 -9.630 0.330 ;
    RECT -11.250 0.000 -11.070 2.095 ;
    RECT -11.250 -0.330 -10.350 0.330 ;
    RECT -11.970 0.000 -11.790 2.095 ;
    RECT -11.970 -0.330 -11.070 0.330 ;
    RECT -12.690 0.000 -12.510 2.095 ;
    RECT -12.690 -0.330 -11.790 0.330 ;
    RECT -13.410 0.000 -13.230 2.095 ;
    RECT -13.410 -0.330 -12.510 0.330 ;
    RECT -14.130 0.000 -13.950 2.095 ;
    RECT -14.130 -0.330 -13.230 0.330 ;
    RECT -7.650 -1.595 -7.470 0.000 ;
    RECT -8.370 -1.595 -8.190 0.000 ;
    RECT -8.370 -0.330 -7.470 0.330 ;
    RECT -9.090 -1.595 -8.910 0.000 ;
    RECT -9.090 -0.330 -8.190 0.330 ;
    RECT -9.810 -1.595 -9.630 0.000 ;
    RECT -9.810 -0.330 -8.910 0.330 ;
    RECT -10.530 -1.595 -10.350 0.000 ;
    RECT -10.530 -0.330 -9.630 0.330 ;
    RECT -11.250 -1.595 -11.070 0.000 ;
    RECT -11.250 -0.330 -10.350 0.330 ;
    RECT -11.970 -1.595 -11.790 0.000 ;
    RECT -11.970 -0.330 -11.070 0.330 ;
    RECT -12.690 -1.595 -12.510 0.000 ;
    RECT -12.690 -0.330 -11.790 0.330 ;
    RECT -13.410 -1.595 -13.230 0.000 ;
    RECT -13.410 -0.330 -12.510 0.330 ;
    RECT -14.130 -1.595 -13.950 0.000 ;
    RECT -14.130 -0.330 -13.230 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT -7.940 -0.130 -7.520 0.290 ;
    LAYER METAL1 ;
    RECT -14.760 2.370 8.280 3.170 ;
    RECT -14.760 -2.670 8.280 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT -8.085 -0.100 -7.615 0.335 ;
    RECT 7.735 -0.010 8.115 0.270 ;
    RECT 1.325 0.000 1.555 0.795 ;
    RECT 0.605 0.565 1.555 0.795 ;
    RECT 1.325 -0.115 8.035 0.115 ;
    RECT -1.555 1.900 0.115 2.130 ;
    RECT -2.995 1.900 -1.325 2.130 ;
    RECT -4.435 1.900 -2.765 2.130 ;
    RECT -5.875 1.900 -4.205 2.130 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT -0.115 1.150 0.115 2.130 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT 1.325 1.150 1.555 2.770 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 0.565 -0.605 1.150 ;
    RECT 2.045 0.000 2.275 1.150 ;
    RECT -0.835 0.565 0.835 0.795 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT -1.555 1.150 -1.325 2.130 ;
    RECT -1.555 1.900 0.115 2.130 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT 2.765 1.150 2.995 2.770 ;
    RECT -2.330 1.035 -1.990 1.265 ;
    RECT 3.430 1.035 3.770 1.265 ;
    RECT -2.275 0.565 -2.045 1.150 ;
    RECT 3.485 0.000 3.715 1.150 ;
    RECT -2.275 0.565 -0.605 0.795 ;
    RECT -3.050 1.035 -2.710 1.265 ;
    RECT -2.995 1.150 -2.765 2.130 ;
    RECT -2.995 1.900 -1.325 2.130 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT 4.205 1.150 4.435 2.770 ;
    RECT -3.770 1.035 -3.430 1.265 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT -3.715 0.565 -3.485 1.150 ;
    RECT 4.925 0.000 5.155 1.150 ;
    RECT -3.715 0.565 -2.045 0.795 ;
    RECT -4.490 1.035 -4.150 1.265 ;
    RECT -4.435 1.150 -4.205 2.130 ;
    RECT -4.435 1.900 -2.765 2.130 ;
    RECT 5.590 1.035 5.930 1.265 ;
    RECT 5.645 1.150 5.875 2.770 ;
    RECT -5.210 1.035 -4.870 1.265 ;
    RECT 6.310 1.035 6.650 1.265 ;
    RECT -5.155 0.565 -4.925 1.150 ;
    RECT 6.365 0.000 6.595 1.150 ;
    RECT -5.155 0.565 -3.485 0.795 ;
    RECT -5.930 1.035 -5.590 1.265 ;
    RECT -5.875 1.150 -5.645 2.130 ;
    RECT -5.875 1.900 -4.205 2.130 ;
    RECT 7.030 1.035 7.370 1.265 ;
    RECT 7.085 1.150 7.315 2.770 ;
    RECT -6.650 1.035 -6.310 1.265 ;
    RECT 7.750 1.035 8.090 1.265 ;
    RECT -6.595 0.565 -6.365 1.150 ;
    RECT 7.805 0.000 8.035 1.150 ;
    RECT -6.595 0.565 -4.925 0.795 ;
    RECT -7.370 1.035 -7.030 1.265 ;
    RECT -7.315 0.565 -7.085 1.150 ;
    RECT -7.315 1.150 -7.085 2.130 ;
    RECT -7.315 1.900 -5.645 2.130 ;
    RECT -8.035 1.150 -7.805 2.770 ;
    RECT -8.090 1.035 -7.750 1.265 ;
    RECT -8.810 1.035 -8.470 1.265 ;
    RECT -8.755 0.565 -8.525 1.150 ;
    RECT -8.755 0.565 -7.085 0.795 ;
    RECT -9.475 1.150 -9.245 2.770 ;
    RECT -9.530 1.035 -9.190 1.265 ;
    RECT -10.250 1.035 -9.910 1.265 ;
    RECT -10.195 0.565 -9.965 1.150 ;
    RECT -10.195 0.565 -8.525 0.795 ;
    RECT -10.915 1.150 -10.685 2.770 ;
    RECT -10.970 1.035 -10.630 1.265 ;
    RECT -11.690 1.035 -11.350 1.265 ;
    RECT -11.635 0.565 -11.405 1.150 ;
    RECT -11.635 0.565 -9.965 0.795 ;
    RECT -12.355 1.150 -12.125 2.770 ;
    RECT -12.410 1.035 -12.070 1.265 ;
    RECT -13.130 1.035 -12.790 1.265 ;
    RECT -13.075 0.565 -12.845 1.150 ;
    RECT -13.075 0.565 -11.405 0.795 ;
    RECT -13.795 1.150 -13.565 2.770 ;
    RECT -13.850 1.035 -13.510 1.265 ;
    RECT -14.570 1.035 -14.230 1.265 ;
    RECT -14.515 0.565 -14.285 1.150 ;
    RECT -14.515 0.565 -12.845 0.795 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT -3.715 -0.560 -2.045 -0.330 ;
    RECT -5.155 -0.560 -3.485 -0.330 ;
    RECT -6.595 -0.560 -4.925 -0.330 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -1.630 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -2.270 0.115 -0.905 ;
    RECT 1.325 -0.905 1.555 0.000 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -0.905 -0.605 -0.330 ;
    RECT 2.045 -1.630 2.275 -0.905 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -1.630 2.275 -1.400 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -2.270 -1.325 -0.905 ;
    RECT 2.765 -0.905 2.995 0.000 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -2.275 -0.905 -2.045 -0.330 ;
    RECT 3.485 -1.630 3.715 -0.905 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT 2.045 -1.630 3.715 -1.400 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -2.270 -2.765 -0.905 ;
    RECT 4.205 -0.905 4.435 0.000 ;
    RECT -3.770 -1.020 -3.430 -0.790 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT -3.715 -0.905 -3.485 -0.330 ;
    RECT 4.925 -1.630 5.155 -0.905 ;
    RECT -3.715 -0.560 -2.045 -0.330 ;
    RECT 3.485 -1.630 5.155 -1.400 ;
    RECT -4.490 -1.020 -4.150 -0.790 ;
    RECT 5.590 -1.020 5.930 -0.790 ;
    RECT -4.435 -2.270 -4.205 -0.905 ;
    RECT 5.645 -0.905 5.875 0.000 ;
    RECT -5.210 -1.020 -4.870 -0.790 ;
    RECT 6.310 -1.020 6.650 -0.790 ;
    RECT -5.155 -0.905 -4.925 -0.330 ;
    RECT 6.365 -1.630 6.595 -0.905 ;
    RECT -5.155 -0.560 -3.485 -0.330 ;
    RECT 4.925 -1.630 6.595 -1.400 ;
    RECT -5.930 -1.020 -5.590 -0.790 ;
    RECT 7.030 -1.020 7.370 -0.790 ;
    RECT -5.875 -2.270 -5.645 -0.905 ;
    RECT 7.085 -0.905 7.315 0.000 ;
    RECT -6.650 -1.020 -6.310 -0.790 ;
    RECT 7.750 -1.020 8.090 -0.790 ;
    RECT -6.595 -0.905 -6.365 -0.330 ;
    RECT 7.805 -1.630 8.035 -0.905 ;
    RECT -6.595 -0.560 -4.925 -0.330 ;
    RECT 6.365 -1.630 8.035 -1.400 ;
    RECT -7.370 -1.020 -7.030 -0.790 ;
    RECT -7.315 -0.905 -7.085 -0.330 ;
    RECT -7.315 -0.560 -5.645 -0.330 ;
    RECT -8.090 -1.020 -7.750 -0.790 ;
    RECT -8.035 -2.270 -7.805 -0.905 ;
    RECT -8.810 -1.020 -8.470 -0.790 ;
    RECT -8.755 -0.905 -8.525 -0.330 ;
    RECT -8.755 -0.560 -7.085 -0.330 ;
    RECT -9.530 -1.020 -9.190 -0.790 ;
    RECT -9.475 -2.270 -9.245 -0.905 ;
    RECT -10.250 -1.020 -9.910 -0.790 ;
    RECT -10.195 -0.905 -9.965 -0.330 ;
    RECT -10.195 -0.560 -8.525 -0.330 ;
    RECT -10.970 -1.020 -10.630 -0.790 ;
    RECT -10.915 -2.270 -10.685 -0.905 ;
    RECT -11.690 -1.020 -11.350 -0.790 ;
    RECT -11.635 -0.905 -11.405 -0.330 ;
    RECT -11.635 -0.560 -9.965 -0.330 ;
    RECT -12.410 -1.020 -12.070 -0.790 ;
    RECT -12.355 -2.270 -12.125 -0.905 ;
    RECT -13.130 -1.020 -12.790 -0.790 ;
    RECT -13.075 -0.905 -12.845 -0.330 ;
    RECT -13.075 -0.560 -11.405 -0.330 ;
    RECT -13.850 -1.020 -13.510 -0.790 ;
    RECT -13.795 -2.270 -13.565 -0.905 ;
    RECT -14.570 -1.020 -14.230 -0.790 ;
    RECT -14.515 -0.905 -14.285 -0.330 ;
    RECT -14.515 -0.560 -12.845 -0.330 ;
    LAYER METAL2 ;
    RECT 7.780 -0.060 8.065 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT -8.085 -0.010 -7.705 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT -7.840 -0.030 -7.620 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT -3.710 2.425 -3.490 2.645 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT -3.710 -2.145 -3.490 -1.925 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT -4.430 2.425 -4.210 2.645 ;
    RECT 5.650 2.425 5.870 2.645 ;
    RECT -4.430 -2.145 -4.210 -1.925 ;
    RECT 5.650 -2.145 5.870 -1.925 ;
    RECT -5.150 2.425 -4.930 2.645 ;
    RECT 6.370 2.425 6.590 2.645 ;
    RECT -5.150 -2.145 -4.930 -1.925 ;
    RECT 6.370 -2.145 6.590 -1.925 ;
    RECT -5.870 2.425 -5.650 2.645 ;
    RECT 7.090 2.425 7.310 2.645 ;
    RECT -5.870 -2.145 -5.650 -1.925 ;
    RECT 7.090 -2.145 7.310 -1.925 ;
    RECT -6.590 2.425 -6.370 2.645 ;
    RECT 7.810 2.425 8.030 2.645 ;
    RECT -6.590 -2.145 -6.370 -1.925 ;
    RECT 7.810 -2.145 8.030 -1.925 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT -2.270 1.040 -2.050 1.260 ;
    RECT 3.490 1.040 3.710 1.260 ;
    RECT -2.990 1.040 -2.770 1.260 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT -3.710 1.040 -3.490 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    RECT -4.430 1.040 -4.210 1.260 ;
    RECT 5.650 1.040 5.870 1.260 ;
    RECT -5.150 1.040 -4.930 1.260 ;
    RECT 6.370 1.040 6.590 1.260 ;
    RECT -5.870 1.040 -5.650 1.260 ;
    RECT 7.090 1.040 7.310 1.260 ;
    RECT -6.590 1.040 -6.370 1.260 ;
    RECT 7.810 1.040 8.030 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT -3.710 -1.015 -3.490 -0.795 ;
    RECT 4.930 -1.015 5.150 -0.795 ;
    RECT -4.430 -1.015 -4.210 -0.795 ;
    RECT 5.650 -1.015 5.870 -0.795 ;
    RECT -5.150 -1.015 -4.930 -0.795 ;
    RECT 6.370 -1.015 6.590 -0.795 ;
    RECT -5.870 -1.015 -5.650 -0.795 ;
    RECT 7.090 -1.015 7.310 -0.795 ;
    RECT -6.590 -1.015 -6.370 -0.795 ;
    RECT 7.810 -1.015 8.030 -0.795 ;
    RECT -7.310 2.425 -7.090 2.645 ;
    RECT -7.310 -2.145 -7.090 -1.925 ;
    RECT -8.030 2.425 -7.810 2.645 ;
    RECT -8.030 -2.145 -7.810 -1.925 ;
    RECT -8.750 2.425 -8.530 2.645 ;
    RECT -8.750 -2.145 -8.530 -1.925 ;
    RECT -9.470 2.425 -9.250 2.645 ;
    RECT -9.470 -2.145 -9.250 -1.925 ;
    RECT -10.190 2.425 -9.970 2.645 ;
    RECT -10.190 -2.145 -9.970 -1.925 ;
    RECT -10.910 2.425 -10.690 2.645 ;
    RECT -10.910 -2.145 -10.690 -1.925 ;
    RECT -11.630 2.425 -11.410 2.645 ;
    RECT -11.630 -2.145 -11.410 -1.925 ;
    RECT -12.350 2.425 -12.130 2.645 ;
    RECT -12.350 -2.145 -12.130 -1.925 ;
    RECT -13.070 2.425 -12.850 2.645 ;
    RECT -13.070 -2.145 -12.850 -1.925 ;
    RECT -13.790 2.425 -13.570 2.645 ;
    RECT -13.790 -2.145 -13.570 -1.925 ;
    RECT -14.510 2.425 -14.290 2.645 ;
    RECT -14.510 -2.145 -14.290 -1.925 ;
    RECT -7.310 1.040 -7.090 1.260 ;
    RECT -8.030 1.040 -7.810 1.260 ;
    RECT -8.750 1.040 -8.530 1.260 ;
    RECT -9.470 1.040 -9.250 1.260 ;
    RECT -10.190 1.040 -9.970 1.260 ;
    RECT -10.910 1.040 -10.690 1.260 ;
    RECT -11.630 1.040 -11.410 1.260 ;
    RECT -12.350 1.040 -12.130 1.260 ;
    RECT -13.070 1.040 -12.850 1.260 ;
    RECT -13.790 1.040 -13.570 1.260 ;
    RECT -14.510 1.040 -14.290 1.260 ;
    RECT -7.310 -1.015 -7.090 -0.795 ;
    RECT -8.030 -1.015 -7.810 -0.795 ;
    RECT -8.750 -1.015 -8.530 -0.795 ;
    RECT -9.470 -1.015 -9.250 -0.795 ;
    RECT -10.190 -1.015 -9.970 -0.795 ;
    RECT -10.910 -1.015 -10.690 -0.795 ;
    RECT -11.630 -1.015 -11.410 -0.795 ;
    RECT -12.350 -1.015 -12.130 -0.795 ;
    RECT -13.070 -1.015 -12.850 -0.795 ;
    RECT -13.790 -1.015 -13.570 -0.795 ;
    RECT -14.510 -1.015 -14.290 -0.795 ;
    LAYER VIA12 ;
    RECT 7.795 0.000 8.055 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT -8.025 0.000 -7.765 0.260 ;
  END
END oai21_1
MACRO oai22_1
  CLASS CORE ;
  FOREIGN oai22_1 -14.760 -2.270 ;
  ORIGIN 14.760 2.270 ;
  SIZE 30.960 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -14.760 2.370 16.200 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -14.760 -2.670 16.200 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 15.700 -0.060 15.985 0.320 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    END
  END in0
  PIN in1
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -8.085 -0.010 -7.705 0.270 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    END
  END in2
  PIN in3
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT 8.475 -0.010 8.855 0.270 ;
    END
  END in3
  OBS
    LAYER NWELL ;
    RECT -15.480 0.000 16.920 3.310 ;
    LAYER NIMP ;
    RECT -14.790 -1.725 16.230 0.000 ;
    RECT -14.860 2.225 16.300 2.990 ;
    LAYER PIMP ;
    RECT -14.790 0.000 16.230 2.225 ;
    RECT -14.860 -2.490 16.300 -1.725 ;
    LAYER N2V ;
    RECT -14.790 -1.725 16.230 0.000 ;
    LAYER P2V ;
    RECT -14.790 0.000 16.230 2.225 ;
    LAYER DIFF ;
    RECT -14.760 -2.380 16.200 -1.825 ;
    RECT -6.690 0.430 8.130 1.875 ;
    RECT 8.430 0.430 16.050 1.875 ;
    RECT -14.610 0.430 -6.990 1.875 ;
    RECT -14.760 2.325 16.200 2.880 ;
    RECT -14.610 -1.375 16.050 -0.430 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.095 ;
    RECT 0.990 0.000 1.170 2.095 ;
    RECT -0.450 0.000 -0.270 2.095 ;
    RECT 1.710 0.000 1.890 2.095 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 0.000 -0.990 2.095 ;
    RECT 2.430 0.000 2.610 2.095 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 0.000 -1.710 2.095 ;
    RECT 3.150 0.000 3.330 2.095 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 0.000 -2.430 2.095 ;
    RECT 3.870 0.000 4.050 2.095 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 0.000 -3.150 2.095 ;
    RECT 4.590 0.000 4.770 2.095 ;
    RECT -3.330 -0.330 -2.430 0.330 ;
    RECT 3.870 -0.330 4.770 0.330 ;
    RECT -4.050 0.000 -3.870 2.095 ;
    RECT 5.310 0.000 5.490 2.095 ;
    RECT -4.050 -0.330 -3.150 0.330 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT -4.770 0.000 -4.590 2.095 ;
    RECT 6.030 0.000 6.210 2.095 ;
    RECT -4.770 -0.330 -3.870 0.330 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT -5.490 0.000 -5.310 2.095 ;
    RECT 6.750 0.000 6.930 2.095 ;
    RECT -5.490 -0.330 -4.590 0.330 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT -6.210 0.000 -6.030 2.095 ;
    RECT 7.470 0.000 7.650 2.095 ;
    RECT -6.210 -0.330 -5.310 0.330 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT 0.270 -1.595 0.450 0.000 ;
    RECT 0.990 -1.595 1.170 0.000 ;
    RECT -0.450 -1.595 -0.270 0.000 ;
    RECT 1.710 -1.595 1.890 0.000 ;
    RECT -0.450 -0.330 0.450 0.330 ;
    RECT 0.990 -0.330 1.890 0.330 ;
    RECT -1.170 -1.595 -0.990 0.000 ;
    RECT 2.430 -1.595 2.610 0.000 ;
    RECT -1.170 -0.330 -0.270 0.330 ;
    RECT 1.710 -0.330 2.610 0.330 ;
    RECT -1.890 -1.595 -1.710 0.000 ;
    RECT 3.150 -1.595 3.330 0.000 ;
    RECT -1.890 -0.330 -0.990 0.330 ;
    RECT 2.430 -0.330 3.330 0.330 ;
    RECT -2.610 -1.595 -2.430 0.000 ;
    RECT 3.870 -1.595 4.050 0.000 ;
    RECT -2.610 -0.330 -1.710 0.330 ;
    RECT 3.150 -0.330 4.050 0.330 ;
    RECT -3.330 -1.595 -3.150 0.000 ;
    RECT 4.590 -1.595 4.770 0.000 ;
    RECT -3.330 -0.330 -2.430 0.330 ;
    RECT 3.870 -0.330 4.770 0.330 ;
    RECT -4.050 -1.595 -3.870 0.000 ;
    RECT 5.310 -1.595 5.490 0.000 ;
    RECT -4.050 -0.330 -3.150 0.330 ;
    RECT 4.590 -0.330 5.490 0.330 ;
    RECT -4.770 -1.595 -4.590 0.000 ;
    RECT 6.030 -1.595 6.210 0.000 ;
    RECT -4.770 -0.330 -3.870 0.330 ;
    RECT 5.310 -0.330 6.210 0.330 ;
    RECT -5.490 -1.595 -5.310 0.000 ;
    RECT 6.750 -1.595 6.930 0.000 ;
    RECT -5.490 -0.330 -4.590 0.330 ;
    RECT 6.030 -0.330 6.930 0.330 ;
    RECT -6.210 -1.595 -6.030 0.000 ;
    RECT 7.470 -1.595 7.650 0.000 ;
    RECT -6.210 -0.330 -5.310 0.330 ;
    RECT 6.750 -0.330 7.650 0.330 ;
    RECT -7.650 0.000 -7.470 2.095 ;
    RECT 8.910 0.000 9.090 2.095 ;
    RECT -8.370 0.000 -8.190 2.095 ;
    RECT 9.630 0.000 9.810 2.095 ;
    RECT -8.370 -0.330 -7.470 0.330 ;
    RECT 8.910 -0.330 9.810 0.330 ;
    RECT -9.090 0.000 -8.910 2.095 ;
    RECT 10.350 0.000 10.530 2.095 ;
    RECT -9.090 -0.330 -8.190 0.330 ;
    RECT 9.630 -0.330 10.530 0.330 ;
    RECT -9.810 0.000 -9.630 2.095 ;
    RECT 11.070 0.000 11.250 2.095 ;
    RECT -9.810 -0.330 -8.910 0.330 ;
    RECT 10.350 -0.330 11.250 0.330 ;
    RECT -10.530 0.000 -10.350 2.095 ;
    RECT 11.790 0.000 11.970 2.095 ;
    RECT -10.530 -0.330 -9.630 0.330 ;
    RECT 11.070 -0.330 11.970 0.330 ;
    RECT -11.250 0.000 -11.070 2.095 ;
    RECT 12.510 0.000 12.690 2.095 ;
    RECT -11.250 -0.330 -10.350 0.330 ;
    RECT 11.790 -0.330 12.690 0.330 ;
    RECT -11.970 0.000 -11.790 2.095 ;
    RECT 13.230 0.000 13.410 2.095 ;
    RECT -11.970 -0.330 -11.070 0.330 ;
    RECT 12.510 -0.330 13.410 0.330 ;
    RECT -12.690 0.000 -12.510 2.095 ;
    RECT 13.950 0.000 14.130 2.095 ;
    RECT -12.690 -0.330 -11.790 0.330 ;
    RECT 13.230 -0.330 14.130 0.330 ;
    RECT -13.410 0.000 -13.230 2.095 ;
    RECT 14.670 0.000 14.850 2.095 ;
    RECT -13.410 -0.330 -12.510 0.330 ;
    RECT 13.950 -0.330 14.850 0.330 ;
    RECT -14.130 0.000 -13.950 2.095 ;
    RECT 15.390 0.000 15.570 2.095 ;
    RECT -14.130 -0.330 -13.230 0.330 ;
    RECT 14.670 -0.330 15.570 0.330 ;
    RECT -7.650 -1.595 -7.470 0.000 ;
    RECT 8.910 -1.595 9.090 0.000 ;
    RECT -8.370 -1.595 -8.190 0.000 ;
    RECT 9.630 -1.595 9.810 0.000 ;
    RECT -8.370 -0.330 -7.470 0.330 ;
    RECT 8.910 -0.330 9.810 0.330 ;
    RECT -9.090 -1.595 -8.910 0.000 ;
    RECT 10.350 -1.595 10.530 0.000 ;
    RECT -9.090 -0.330 -8.190 0.330 ;
    RECT 9.630 -0.330 10.530 0.330 ;
    RECT -9.810 -1.595 -9.630 0.000 ;
    RECT 11.070 -1.595 11.250 0.000 ;
    RECT -9.810 -0.330 -8.910 0.330 ;
    RECT 10.350 -0.330 11.250 0.330 ;
    RECT -10.530 -1.595 -10.350 0.000 ;
    RECT 11.790 -1.595 11.970 0.000 ;
    RECT -10.530 -0.330 -9.630 0.330 ;
    RECT 11.070 -0.330 11.970 0.330 ;
    RECT -11.250 -1.595 -11.070 0.000 ;
    RECT 12.510 -1.595 12.690 0.000 ;
    RECT -11.250 -0.330 -10.350 0.330 ;
    RECT 11.790 -0.330 12.690 0.330 ;
    RECT -11.970 -1.595 -11.790 0.000 ;
    RECT 13.230 -1.595 13.410 0.000 ;
    RECT -11.970 -0.330 -11.070 0.330 ;
    RECT 12.510 -0.330 13.410 0.330 ;
    RECT -12.690 -1.595 -12.510 0.000 ;
    RECT 13.950 -1.595 14.130 0.000 ;
    RECT -12.690 -0.330 -11.790 0.330 ;
    RECT 13.230 -0.330 14.130 0.330 ;
    RECT -13.410 -1.595 -13.230 0.000 ;
    RECT 14.670 -1.595 14.850 0.000 ;
    RECT -13.410 -0.330 -12.510 0.330 ;
    RECT 13.950 -0.330 14.850 0.330 ;
    RECT -14.130 -1.595 -13.950 0.000 ;
    RECT 15.390 -1.595 15.570 0.000 ;
    RECT -14.130 -0.330 -13.230 0.330 ;
    RECT 14.670 -0.330 15.570 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    RECT 0.700 -0.130 1.120 0.290 ;
    RECT 8.620 -0.130 9.040 0.290 ;
    RECT -7.940 -0.130 -7.520 0.290 ;
    LAYER METAL1 ;
    RECT -14.760 2.370 16.200 3.170 ;
    RECT -14.760 -2.670 16.200 -1.870 ;
    RECT -0.165 -0.100 0.305 0.335 ;
    RECT 0.555 -0.100 1.025 0.335 ;
    RECT 8.475 -0.100 8.945 0.335 ;
    RECT -8.085 -0.100 -7.615 0.335 ;
    RECT 15.655 -0.010 16.035 0.270 ;
    RECT 15.725 -0.560 15.955 0.000 ;
    RECT 1.325 -0.560 15.955 -0.330 ;
    RECT 7.085 -0.560 7.315 0.795 ;
    RECT -0.115 1.900 1.555 2.130 ;
    RECT -0.115 1.900 1.555 2.130 ;
    RECT -1.555 1.900 0.115 2.130 ;
    RECT 1.325 1.900 2.995 2.130 ;
    RECT -2.995 1.900 -1.325 2.130 ;
    RECT 2.765 1.900 4.435 2.130 ;
    RECT -4.435 1.900 -2.765 2.130 ;
    RECT 4.205 1.900 5.875 2.130 ;
    RECT -5.875 1.900 -4.205 2.130 ;
    RECT 5.645 1.900 7.315 2.130 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT 0.605 0.565 0.835 1.150 ;
    RECT 0.605 0.565 2.275 0.795 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT -0.115 1.150 0.115 2.130 ;
    RECT 1.325 1.150 1.555 2.130 ;
    RECT -0.115 1.900 1.555 2.130 ;
    RECT -0.115 1.900 1.555 2.130 ;
    RECT -0.890 1.035 -0.550 1.265 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT -0.835 0.565 -0.605 1.150 ;
    RECT 2.045 0.565 2.275 1.150 ;
    RECT -0.835 0.565 0.835 0.795 ;
    RECT 0.605 0.565 2.275 0.795 ;
    RECT -1.610 1.035 -1.270 1.265 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT -1.555 1.150 -1.325 2.130 ;
    RECT 2.765 1.150 2.995 2.130 ;
    RECT -1.555 1.900 0.115 2.130 ;
    RECT 1.325 1.900 2.995 2.130 ;
    RECT -2.330 1.035 -1.990 1.265 ;
    RECT 3.430 1.035 3.770 1.265 ;
    RECT -2.275 0.565 -2.045 1.150 ;
    RECT 3.485 0.565 3.715 1.150 ;
    RECT -2.275 0.565 -0.605 0.795 ;
    RECT 2.045 0.565 3.715 0.795 ;
    RECT -3.050 1.035 -2.710 1.265 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT -2.995 1.150 -2.765 2.130 ;
    RECT 4.205 1.150 4.435 2.130 ;
    RECT -2.995 1.900 -1.325 2.130 ;
    RECT 2.765 1.900 4.435 2.130 ;
    RECT -3.770 1.035 -3.430 1.265 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT -3.715 0.565 -3.485 1.150 ;
    RECT 4.925 0.565 5.155 1.150 ;
    RECT -3.715 0.565 -2.045 0.795 ;
    RECT 3.485 0.565 5.155 0.795 ;
    RECT -4.490 1.035 -4.150 1.265 ;
    RECT 5.590 1.035 5.930 1.265 ;
    RECT -4.435 1.150 -4.205 2.130 ;
    RECT 5.645 1.150 5.875 2.130 ;
    RECT -4.435 1.900 -2.765 2.130 ;
    RECT 4.205 1.900 5.875 2.130 ;
    RECT -5.210 1.035 -4.870 1.265 ;
    RECT 6.310 1.035 6.650 1.265 ;
    RECT -5.155 0.565 -4.925 1.150 ;
    RECT 6.365 0.565 6.595 1.150 ;
    RECT -5.155 0.565 -3.485 0.795 ;
    RECT 4.925 0.565 6.595 0.795 ;
    RECT -5.930 1.035 -5.590 1.265 ;
    RECT 7.030 1.035 7.370 1.265 ;
    RECT -5.875 1.150 -5.645 2.130 ;
    RECT 7.085 1.150 7.315 2.130 ;
    RECT -5.875 1.900 -4.205 2.130 ;
    RECT 5.645 1.900 7.315 2.130 ;
    RECT -6.650 1.035 -6.310 1.265 ;
    RECT 7.750 1.035 8.090 1.265 ;
    RECT -6.595 0.565 -6.365 1.150 ;
    RECT 7.805 0.565 8.035 1.150 ;
    RECT -6.595 0.565 -4.925 0.795 ;
    RECT 6.365 0.565 8.035 0.795 ;
    RECT -7.370 1.035 -7.030 1.265 ;
    RECT 8.470 1.035 8.810 1.265 ;
    RECT -7.315 0.565 -7.085 1.150 ;
    RECT 8.525 0.565 8.755 1.150 ;
    RECT -7.315 1.150 -7.085 2.130 ;
    RECT 8.525 1.150 8.755 2.130 ;
    RECT -7.315 1.900 -5.645 2.130 ;
    RECT 7.085 1.900 8.755 2.130 ;
    RECT -8.035 1.150 -7.805 2.770 ;
    RECT 9.245 1.150 9.475 2.770 ;
    RECT -8.090 1.035 -7.750 1.265 ;
    RECT 9.190 1.035 9.530 1.265 ;
    RECT -8.810 1.035 -8.470 1.265 ;
    RECT 9.910 1.035 10.250 1.265 ;
    RECT -8.755 0.565 -8.525 1.150 ;
    RECT 9.965 0.565 10.195 1.150 ;
    RECT -8.755 0.565 -7.085 0.795 ;
    RECT 8.525 0.565 10.195 0.795 ;
    RECT -9.475 1.150 -9.245 2.770 ;
    RECT 10.685 1.150 10.915 2.770 ;
    RECT -9.530 1.035 -9.190 1.265 ;
    RECT 10.630 1.035 10.970 1.265 ;
    RECT -10.250 1.035 -9.910 1.265 ;
    RECT 11.350 1.035 11.690 1.265 ;
    RECT -10.195 0.565 -9.965 1.150 ;
    RECT 11.405 0.565 11.635 1.150 ;
    RECT -10.195 0.565 -8.525 0.795 ;
    RECT 9.965 0.565 11.635 0.795 ;
    RECT -10.915 1.150 -10.685 2.770 ;
    RECT 12.125 1.150 12.355 2.770 ;
    RECT -10.970 1.035 -10.630 1.265 ;
    RECT 12.070 1.035 12.410 1.265 ;
    RECT -11.690 1.035 -11.350 1.265 ;
    RECT 12.790 1.035 13.130 1.265 ;
    RECT -11.635 0.565 -11.405 1.150 ;
    RECT 12.845 0.565 13.075 1.150 ;
    RECT -11.635 0.565 -9.965 0.795 ;
    RECT 11.405 0.565 13.075 0.795 ;
    RECT -12.355 1.150 -12.125 2.770 ;
    RECT 13.565 1.150 13.795 2.770 ;
    RECT -12.410 1.035 -12.070 1.265 ;
    RECT 13.510 1.035 13.850 1.265 ;
    RECT -13.130 1.035 -12.790 1.265 ;
    RECT 14.230 1.035 14.570 1.265 ;
    RECT -13.075 0.565 -12.845 1.150 ;
    RECT 14.285 0.565 14.515 1.150 ;
    RECT -13.075 0.565 -11.405 0.795 ;
    RECT 12.845 0.565 14.515 0.795 ;
    RECT -13.795 1.150 -13.565 2.770 ;
    RECT 15.005 1.150 15.235 2.770 ;
    RECT -13.850 1.035 -13.510 1.265 ;
    RECT 14.950 1.035 15.290 1.265 ;
    RECT -14.570 1.035 -14.230 1.265 ;
    RECT 15.670 1.035 16.010 1.265 ;
    RECT -14.515 0.565 -14.285 1.150 ;
    RECT 15.725 0.565 15.955 1.150 ;
    RECT -14.515 0.565 -12.845 0.795 ;
    RECT 14.285 0.565 15.955 0.795 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -1.630 2.275 -1.400 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT 2.045 -1.630 3.715 -1.400 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT -3.715 -0.560 -2.045 -0.330 ;
    RECT 3.485 -1.630 5.155 -1.400 ;
    RECT 4.205 -0.560 5.875 -0.330 ;
    RECT -5.155 -0.560 -3.485 -0.330 ;
    RECT 4.925 -1.630 6.595 -1.400 ;
    RECT 5.645 -0.560 7.315 -0.330 ;
    RECT -6.595 -0.560 -4.925 -0.330 ;
    RECT 6.365 -1.630 8.035 -1.400 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 -0.330 ;
    RECT 0.605 -1.630 0.835 -0.905 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT -0.115 -2.270 0.115 -0.905 ;
    RECT 1.325 -0.905 1.555 -0.330 ;
    RECT -0.890 -1.020 -0.550 -0.790 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT -0.835 -0.905 -0.605 -0.330 ;
    RECT 2.045 -1.630 2.275 -0.905 ;
    RECT -0.835 -0.560 0.835 -0.330 ;
    RECT 0.605 -1.630 2.275 -1.400 ;
    RECT -1.610 -1.020 -1.270 -0.790 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT -1.555 -2.270 -1.325 -0.905 ;
    RECT 2.765 -0.905 2.995 -0.330 ;
    RECT 1.325 -0.560 2.995 -0.330 ;
    RECT -2.330 -1.020 -1.990 -0.790 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT -2.275 -0.905 -2.045 -0.330 ;
    RECT 3.485 -1.630 3.715 -0.905 ;
    RECT -2.275 -0.560 -0.605 -0.330 ;
    RECT 2.045 -1.630 3.715 -1.400 ;
    RECT -3.050 -1.020 -2.710 -0.790 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT -2.995 -2.270 -2.765 -0.905 ;
    RECT 4.205 -0.905 4.435 -0.330 ;
    RECT 2.765 -0.560 4.435 -0.330 ;
    RECT -3.770 -1.020 -3.430 -0.790 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT -3.715 -0.905 -3.485 -0.330 ;
    RECT 4.925 -1.630 5.155 -0.905 ;
    RECT -3.715 -0.560 -2.045 -0.330 ;
    RECT 3.485 -1.630 5.155 -1.400 ;
    RECT -4.490 -1.020 -4.150 -0.790 ;
    RECT 5.590 -1.020 5.930 -0.790 ;
    RECT -4.435 -2.270 -4.205 -0.905 ;
    RECT 5.645 -0.905 5.875 -0.330 ;
    RECT 4.205 -0.560 5.875 -0.330 ;
    RECT -5.210 -1.020 -4.870 -0.790 ;
    RECT 6.310 -1.020 6.650 -0.790 ;
    RECT -5.155 -0.905 -4.925 -0.330 ;
    RECT 6.365 -1.630 6.595 -0.905 ;
    RECT -5.155 -0.560 -3.485 -0.330 ;
    RECT 4.925 -1.630 6.595 -1.400 ;
    RECT -5.930 -1.020 -5.590 -0.790 ;
    RECT 7.030 -1.020 7.370 -0.790 ;
    RECT -5.875 -2.270 -5.645 -0.905 ;
    RECT 7.085 -0.905 7.315 -0.330 ;
    RECT 5.645 -0.560 7.315 -0.330 ;
    RECT -6.650 -1.020 -6.310 -0.790 ;
    RECT 7.750 -1.020 8.090 -0.790 ;
    RECT -6.595 -0.905 -6.365 -0.330 ;
    RECT 7.805 -1.630 8.035 -0.905 ;
    RECT -6.595 -0.560 -4.925 -0.330 ;
    RECT 6.365 -1.630 8.035 -1.400 ;
    RECT -7.370 -1.020 -7.030 -0.790 ;
    RECT 8.470 -1.020 8.810 -0.790 ;
    RECT -7.315 -0.905 -7.085 -0.330 ;
    RECT 8.525 -1.630 8.755 -0.905 ;
    RECT -7.315 -0.560 -5.645 -0.330 ;
    RECT 7.085 -1.630 8.755 -1.400 ;
    RECT -8.090 -1.020 -7.750 -0.790 ;
    RECT 9.190 -1.020 9.530 -0.790 ;
    RECT -8.035 -2.270 -7.805 -0.905 ;
    RECT 9.245 -0.905 9.475 -0.330 ;
    RECT 7.085 -0.560 9.475 -0.330 ;
    RECT -8.810 -1.020 -8.470 -0.790 ;
    RECT 9.910 -1.020 10.250 -0.790 ;
    RECT -8.755 -0.905 -8.525 -0.330 ;
    RECT 9.965 -1.630 10.195 -0.905 ;
    RECT -8.755 -0.560 -7.085 -0.330 ;
    RECT 8.525 -1.630 10.195 -1.400 ;
    RECT -9.530 -1.020 -9.190 -0.790 ;
    RECT 10.630 -1.020 10.970 -0.790 ;
    RECT -9.475 -2.270 -9.245 -0.905 ;
    RECT 10.685 -0.905 10.915 -0.330 ;
    RECT 8.525 -0.560 10.915 -0.330 ;
    RECT -10.250 -1.020 -9.910 -0.790 ;
    RECT 11.350 -1.020 11.690 -0.790 ;
    RECT -10.195 -0.905 -9.965 -0.330 ;
    RECT 11.405 -1.630 11.635 -0.905 ;
    RECT -10.195 -0.560 -8.525 -0.330 ;
    RECT 9.965 -1.630 11.635 -1.400 ;
    RECT -10.970 -1.020 -10.630 -0.790 ;
    RECT 12.070 -1.020 12.410 -0.790 ;
    RECT -10.915 -2.270 -10.685 -0.905 ;
    RECT 12.125 -0.905 12.355 -0.330 ;
    RECT 9.965 -0.560 12.355 -0.330 ;
    RECT -11.690 -1.020 -11.350 -0.790 ;
    RECT 12.790 -1.020 13.130 -0.790 ;
    RECT -11.635 -0.905 -11.405 -0.330 ;
    RECT 12.845 -1.630 13.075 -0.905 ;
    RECT -11.635 -0.560 -9.965 -0.330 ;
    RECT 11.405 -1.630 13.075 -1.400 ;
    RECT -12.410 -1.020 -12.070 -0.790 ;
    RECT 13.510 -1.020 13.850 -0.790 ;
    RECT -12.355 -2.270 -12.125 -0.905 ;
    RECT 13.565 -0.905 13.795 -0.330 ;
    RECT 11.405 -0.560 13.795 -0.330 ;
    RECT -13.130 -1.020 -12.790 -0.790 ;
    RECT 14.230 -1.020 14.570 -0.790 ;
    RECT -13.075 -0.905 -12.845 -0.330 ;
    RECT 14.285 -1.630 14.515 -0.905 ;
    RECT -13.075 -0.560 -11.405 -0.330 ;
    RECT 12.845 -1.630 14.515 -1.400 ;
    RECT -13.850 -1.020 -13.510 -0.790 ;
    RECT 14.950 -1.020 15.290 -0.790 ;
    RECT -13.795 -2.270 -13.565 -0.905 ;
    RECT 15.005 -0.905 15.235 -0.330 ;
    RECT 12.845 -0.560 15.235 -0.330 ;
    RECT -14.570 -1.020 -14.230 -0.790 ;
    RECT 15.670 -1.020 16.010 -0.790 ;
    RECT -14.515 -0.905 -14.285 -0.330 ;
    RECT 15.725 -1.630 15.955 -0.905 ;
    RECT -14.515 -0.560 -12.845 -0.330 ;
    RECT 14.285 -1.630 15.955 -1.400 ;
    LAYER METAL2 ;
    RECT 15.700 -0.060 15.985 0.320 ;
    RECT -0.165 -0.010 0.215 0.270 ;
    RECT 0.555 -0.010 0.935 0.270 ;
    RECT 8.475 -0.010 8.855 0.270 ;
    RECT -8.085 -0.010 -7.705 0.270 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT 0.800 -0.030 1.020 0.190 ;
    RECT 8.720 -0.030 8.940 0.190 ;
    RECT -7.840 -0.030 -7.620 0.190 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT -0.830 2.425 -0.610 2.645 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT -0.830 -2.145 -0.610 -1.925 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT -1.550 2.425 -1.330 2.645 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT -1.550 -2.145 -1.330 -1.925 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT -2.270 2.425 -2.050 2.645 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT -2.270 -2.145 -2.050 -1.925 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT -2.990 2.425 -2.770 2.645 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT -2.990 -2.145 -2.770 -1.925 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT -3.710 2.425 -3.490 2.645 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT -3.710 -2.145 -3.490 -1.925 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT -4.430 2.425 -4.210 2.645 ;
    RECT 5.650 2.425 5.870 2.645 ;
    RECT -4.430 -2.145 -4.210 -1.925 ;
    RECT 5.650 -2.145 5.870 -1.925 ;
    RECT -5.150 2.425 -4.930 2.645 ;
    RECT 6.370 2.425 6.590 2.645 ;
    RECT -5.150 -2.145 -4.930 -1.925 ;
    RECT 6.370 -2.145 6.590 -1.925 ;
    RECT -5.870 2.425 -5.650 2.645 ;
    RECT 7.090 2.425 7.310 2.645 ;
    RECT -5.870 -2.145 -5.650 -1.925 ;
    RECT 7.090 -2.145 7.310 -1.925 ;
    RECT -6.590 2.425 -6.370 2.645 ;
    RECT 7.810 2.425 8.030 2.645 ;
    RECT -6.590 -2.145 -6.370 -1.925 ;
    RECT 7.810 -2.145 8.030 -1.925 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT -0.830 1.040 -0.610 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT -1.550 1.040 -1.330 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT -2.270 1.040 -2.050 1.260 ;
    RECT 3.490 1.040 3.710 1.260 ;
    RECT -2.990 1.040 -2.770 1.260 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT -3.710 1.040 -3.490 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    RECT -4.430 1.040 -4.210 1.260 ;
    RECT 5.650 1.040 5.870 1.260 ;
    RECT -5.150 1.040 -4.930 1.260 ;
    RECT 6.370 1.040 6.590 1.260 ;
    RECT -5.870 1.040 -5.650 1.260 ;
    RECT 7.090 1.040 7.310 1.260 ;
    RECT -6.590 1.040 -6.370 1.260 ;
    RECT 7.810 1.040 8.030 1.260 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT 0.610 -1.015 0.830 -0.795 ;
    RECT -0.110 -1.015 0.110 -0.795 ;
    RECT 1.330 -1.015 1.550 -0.795 ;
    RECT -0.830 -1.015 -0.610 -0.795 ;
    RECT 2.050 -1.015 2.270 -0.795 ;
    RECT -1.550 -1.015 -1.330 -0.795 ;
    RECT 2.770 -1.015 2.990 -0.795 ;
    RECT -2.270 -1.015 -2.050 -0.795 ;
    RECT 3.490 -1.015 3.710 -0.795 ;
    RECT -2.990 -1.015 -2.770 -0.795 ;
    RECT 4.210 -1.015 4.430 -0.795 ;
    RECT -3.710 -1.015 -3.490 -0.795 ;
    RECT 4.930 -1.015 5.150 -0.795 ;
    RECT -4.430 -1.015 -4.210 -0.795 ;
    RECT 5.650 -1.015 5.870 -0.795 ;
    RECT -5.150 -1.015 -4.930 -0.795 ;
    RECT 6.370 -1.015 6.590 -0.795 ;
    RECT -5.870 -1.015 -5.650 -0.795 ;
    RECT 7.090 -1.015 7.310 -0.795 ;
    RECT -6.590 -1.015 -6.370 -0.795 ;
    RECT 7.810 -1.015 8.030 -0.795 ;
    RECT -7.310 2.425 -7.090 2.645 ;
    RECT 8.530 2.425 8.750 2.645 ;
    RECT -7.310 -2.145 -7.090 -1.925 ;
    RECT 8.530 -2.145 8.750 -1.925 ;
    RECT -8.030 2.425 -7.810 2.645 ;
    RECT 9.250 2.425 9.470 2.645 ;
    RECT -8.030 -2.145 -7.810 -1.925 ;
    RECT 9.250 -2.145 9.470 -1.925 ;
    RECT -8.750 2.425 -8.530 2.645 ;
    RECT 9.970 2.425 10.190 2.645 ;
    RECT -8.750 -2.145 -8.530 -1.925 ;
    RECT 9.970 -2.145 10.190 -1.925 ;
    RECT -9.470 2.425 -9.250 2.645 ;
    RECT 10.690 2.425 10.910 2.645 ;
    RECT -9.470 -2.145 -9.250 -1.925 ;
    RECT 10.690 -2.145 10.910 -1.925 ;
    RECT -10.190 2.425 -9.970 2.645 ;
    RECT 11.410 2.425 11.630 2.645 ;
    RECT -10.190 -2.145 -9.970 -1.925 ;
    RECT 11.410 -2.145 11.630 -1.925 ;
    RECT -10.910 2.425 -10.690 2.645 ;
    RECT 12.130 2.425 12.350 2.645 ;
    RECT -10.910 -2.145 -10.690 -1.925 ;
    RECT 12.130 -2.145 12.350 -1.925 ;
    RECT -11.630 2.425 -11.410 2.645 ;
    RECT 12.850 2.425 13.070 2.645 ;
    RECT -11.630 -2.145 -11.410 -1.925 ;
    RECT 12.850 -2.145 13.070 -1.925 ;
    RECT -12.350 2.425 -12.130 2.645 ;
    RECT 13.570 2.425 13.790 2.645 ;
    RECT -12.350 -2.145 -12.130 -1.925 ;
    RECT 13.570 -2.145 13.790 -1.925 ;
    RECT -13.070 2.425 -12.850 2.645 ;
    RECT 14.290 2.425 14.510 2.645 ;
    RECT -13.070 -2.145 -12.850 -1.925 ;
    RECT 14.290 -2.145 14.510 -1.925 ;
    RECT -13.790 2.425 -13.570 2.645 ;
    RECT 15.010 2.425 15.230 2.645 ;
    RECT -13.790 -2.145 -13.570 -1.925 ;
    RECT 15.010 -2.145 15.230 -1.925 ;
    RECT -14.510 2.425 -14.290 2.645 ;
    RECT 15.730 2.425 15.950 2.645 ;
    RECT -14.510 -2.145 -14.290 -1.925 ;
    RECT 15.730 -2.145 15.950 -1.925 ;
    RECT -7.310 1.040 -7.090 1.260 ;
    RECT 8.530 1.040 8.750 1.260 ;
    RECT -8.030 1.040 -7.810 1.260 ;
    RECT 9.250 1.040 9.470 1.260 ;
    RECT -8.750 1.040 -8.530 1.260 ;
    RECT 9.970 1.040 10.190 1.260 ;
    RECT -9.470 1.040 -9.250 1.260 ;
    RECT 10.690 1.040 10.910 1.260 ;
    RECT -10.190 1.040 -9.970 1.260 ;
    RECT 11.410 1.040 11.630 1.260 ;
    RECT -10.910 1.040 -10.690 1.260 ;
    RECT 12.130 1.040 12.350 1.260 ;
    RECT -11.630 1.040 -11.410 1.260 ;
    RECT 12.850 1.040 13.070 1.260 ;
    RECT -12.350 1.040 -12.130 1.260 ;
    RECT 13.570 1.040 13.790 1.260 ;
    RECT -13.070 1.040 -12.850 1.260 ;
    RECT 14.290 1.040 14.510 1.260 ;
    RECT -13.790 1.040 -13.570 1.260 ;
    RECT 15.010 1.040 15.230 1.260 ;
    RECT -14.510 1.040 -14.290 1.260 ;
    RECT 15.730 1.040 15.950 1.260 ;
    RECT -7.310 -1.015 -7.090 -0.795 ;
    RECT 8.530 -1.015 8.750 -0.795 ;
    RECT -8.030 -1.015 -7.810 -0.795 ;
    RECT 9.250 -1.015 9.470 -0.795 ;
    RECT -8.750 -1.015 -8.530 -0.795 ;
    RECT 9.970 -1.015 10.190 -0.795 ;
    RECT -9.470 -1.015 -9.250 -0.795 ;
    RECT 10.690 -1.015 10.910 -0.795 ;
    RECT -10.190 -1.015 -9.970 -0.795 ;
    RECT 11.410 -1.015 11.630 -0.795 ;
    RECT -10.910 -1.015 -10.690 -0.795 ;
    RECT 12.130 -1.015 12.350 -0.795 ;
    RECT -11.630 -1.015 -11.410 -0.795 ;
    RECT 12.850 -1.015 13.070 -0.795 ;
    RECT -12.350 -1.015 -12.130 -0.795 ;
    RECT 13.570 -1.015 13.790 -0.795 ;
    RECT -13.070 -1.015 -12.850 -0.795 ;
    RECT 14.290 -1.015 14.510 -0.795 ;
    RECT -13.790 -1.015 -13.570 -0.795 ;
    RECT 15.010 -1.015 15.230 -0.795 ;
    RECT -14.510 -1.015 -14.290 -0.795 ;
    RECT 15.730 -1.015 15.950 -0.795 ;
    LAYER VIA12 ;
    RECT 15.715 0.000 15.975 0.260 ;
    RECT -0.105 0.000 0.155 0.260 ;
    RECT 0.615 0.000 0.875 0.260 ;
    RECT 8.535 0.000 8.795 0.260 ;
    RECT -8.025 0.000 -7.765 0.260 ;
  END
END oai22_1
MACRO filler
  CLASS CORE ;
  FOREIGN filler -20.000 -22.000 ;
  ORIGIN 20.000 22.000 ;
  SIZE 16.000 BY 44.000 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -20.000 20.000 -4.000 24.000 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -20.000 -24.000 -4.000 -20.000 ;
    END
  END gnd!
  PIN shield_0
    DIRECTION INOUT ;
    PORT
    LAYER METAL2 ;
    RECT -6.000 -24.000 -2.000 24.000 ;
    END
  END shield_0
  PIN shield_1
    DIRECTION INOUT ;
    PORT
    LAYER METAL2 ;
    RECT -22.000 -24.000 -18.000 24.000 ;
    END
  END shield_1
  OBS
    LAYER NWELL ;
    RECT -24.000 0.000 0.000 28.000 ;
    LAYER NIMP ;
    RECT -20.000 18.000 -4.000 26.000 ;
    RECT -20.000 -18.000 -4.000 0.000 ;
    LAYER PIMP ;
    RECT -20.000 -26.000 -4.000 -18.000 ;
    RECT -20.000 0.000 -4.000 18.000 ;
    LAYER DIFF ;
    RECT -18.000 20.000 -6.000 24.000 ;
    LAYER DIFF ;
    RECT -18.000 -24.000 -6.000 -20.000 ;
    LAYER CONT ;
    RECT -9.000 21.000 -7.000 23.000 ;
    RECT -9.000 -23.000 -7.000 -21.000 ;
    RECT -17.000 21.000 -15.000 23.000 ;
    RECT -17.000 -23.000 -15.000 -21.000 ;
  END
END filler
END LIBRARY
