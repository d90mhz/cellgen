module invload(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_1(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_2(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_3(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_4(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_5(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_6(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_7(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_8(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_9(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_10(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_11(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_12(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_13(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_14(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module inv1x_15(in0, out);
input in0;
output out;
assign out = ~(in0);
endmodule

module nand2_1(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_2(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_3(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_4(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_5(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_6(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_7(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_8(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_9(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_10(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_11(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand2_12(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 & in1);
endmodule

module nand3_1(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_2(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_3(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_4(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_5(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_6(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_7(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_8(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand3_9(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 & in1 & in2);
endmodule

module nand4_1(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~(in0 & in1 & in2 & in3);
endmodule

module nand4_2(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~(in0 & in1 & in2 & in3);
endmodule

module nand4_3(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~(in0 & in1 & in2 & in3);
endmodule

module nand4_4(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~(in0 & in1 & in2 & in3);
endmodule

module nand4_5(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~(in0 & in1 & in2 & in3);
endmodule

module nor2_1(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 | in1);
endmodule

module nor2_2(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 | in1);
endmodule

module nor2_3(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 | in1);
endmodule

module nor2_4(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 | in1);
endmodule

module nor2_5(in0, in1, out);
input in0, in1;
output out;
assign out = ~(in0 | in1);
endmodule

module nor3_1(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 | in1 | in2);
endmodule

module nor3_2(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~(in0 | in1 | in2);
endmodule

module aoi21_1(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_2(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_3(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_4(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_5(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_6(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_7(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_8(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_9(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi21_10(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 & in1) | in2);
endmodule

module aoi22_1(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~((in0 & in1) | (in2 & in3));
endmodule

module oai21_1(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 | in1) & in2);
endmodule

module oai21_2(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 | in1) & in2);
endmodule

module oai21_3(in0, in1, in2, out);
input in0, in1, in2;
output out;
assign out = ~((in0 | in1) & in2);
endmodule

module oai22_1(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~((in0 | in1) & (in2 | in3));
endmodule

module oai22_2(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~((in0 | in1) & (in2 | in3));
endmodule

module oai22_3(in0, in1, in2, in3, out);
input in0, in1, in2, in3;
output out;
assign out = ~((in0 | in1) & (in2 | in3));
endmodule

module too_large ( a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0);
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, q, r, s, t, u, v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0; 
output n0, o0, p0; 

nand2_1 U1 ( .in0(net801), .in1(net934), .out(net820));
nand2_1 U2 ( .in0(net820), .in1(net821), .out(net819));
oai21_1 U3 ( .in0(net931), .in1(net731), .in2(net745), .out(net934));
inv1x_1 U4 ( .in0(net731), .out(net830));
inv1x_2 U5 ( .in0(net741), .out(net931));
inv1x_3 U6 ( .in0(net931), .out(net3006));
nor2_1 U7 ( .in0(net754), .in1(n405), .out(net801));
inv1x_2 U8 ( .in0(n406), .out(n405));
nor2_2 U9 ( .in0(net754), .in1(n405), .out(net825));
nand2_2 U10 ( .in0(net673), .in1(net680), .out(n406));
inv1x_4 U11 ( .in0(d0), .out(net680));
inv1x_5 U12 ( .in0(net723), .out(net754));
nand4_1 U13 ( .in0(net891), .in1(w), .in2(net800), .in3(n407), .out(net745));
nand3_1 U14 ( .in0(net743), .in1(net744), .in2(net745), .out(net742));
nand3_2 U15 ( .in0(net659), .in1(net966), .in2(net981), .out(n407));
inv1x_5 U16 ( .in0(net875), .out(net981));
inv1x_6 U17 ( .in0(net2984), .out(net875));
oai21_1 U18 ( .in0(net873), .in1(net875), .in2(net705), .out(net920));
inv1x_7 U19 ( .in0(net873), .out(net966));
inv1x_8 U20 ( .in0(net733), .out(net873));
nand2_2 U21 ( .in0(net873), .in1(net705), .out(net945));
inv1x_9 U22 ( .in0(net958), .out(net659));
inv1x_10 U23 ( .in0(net1654), .out(net958));
aoi21_1 U24 ( .in0(net958), .in1(net852), .in2(net671), .out(net642));
nand2_3 U25 ( .in0(net958), .in1(net697), .out(net917));
nand3_3 U26 ( .in0(net958), .in1(net926), .in2(net693), .out(net757));
nor2_2 U27 ( .in0(net685), .in1(net680), .out(net800));
inv1x_4 U28 ( .in0(net729), .out(net891));
nand2_4 U29 ( .in0(net1687), .in1(net730), .out(net731));
aoi21_2 U30 ( .in0(net799), .in1(net822), .in2(net819), .out(net646));
nand2_5 U31 ( .in0(v), .in1(net779), .out(net821));
inv1x_2 U32 ( .in0(net821), .out(net783));
inv1x_8 U33 ( .in0(net688), .out(net779));
nand2_6 U34 ( .in0(j0), .in1(net2949), .out(net2984));
aoi21_3 U35 ( .in0(net2956), .in1(net2984), .in2(net2995), .out(net2994));
nand2_4 U36 ( .in0(net2984), .in1(net2956), .out(net2959));
inv1x_9 U37 ( .in0(i0), .out(net2949));
nand2_4 U38 ( .in0(net1592), .in1(net2949), .out(net1636));
nand2_5 U39 ( .in0(net1620), .in1(i0), .out(net733));
inv1x_3 U40 ( .in0(net733), .out(net986));
inv1x_11 U41 ( .in0(y), .out(net1620));
nand2_7 U42 ( .in0(net1655), .in1(net1666), .out(net1654));
nor2_2 U43 ( .in0(net1654), .in1(c0), .out(net684));
inv1x_12 U44 ( .in0(y), .out(net1666));
inv1x_12 U45 ( .in0(a0), .out(net1655));
nand2_5 U46 ( .in0(a0), .in1(net697), .out(net907));
nand2_8 U47 ( .in0(net645), .in1(net646), .out(o0));
nand4_2 U48 ( .in0(net927), .in1(net866), .in2(net928), .in3(n409), .out(net822));
aoi21_3 U49 ( .in0(net797), .in1(net964), .in2(net755), .out(n409));
oai21_1 U50 ( .in0(net693), .in1(net756), .in2(net757), .out(net755));
inv1x_3 U51 ( .in0(u), .out(net693));
nand2_2 U52 ( .in0(net691), .in1(net693), .out(net738));
oai21_2 U53 ( .in0(net693), .in1(net673), .in2(net911), .out(net797));
oai22_1 U54 ( .in0(net680), .in1(net718), .in2(net793), .in3(net794), .out(net926));
nand3_4 U55 ( .in0(l0), .in1(net791), .in2(net795), .out(net794));
nand3_4 U56 ( .in0(net704), .in1(n408), .in2(net652), .out(net793));
inv1x_2 U57 ( .in0(a), .out(n408));
nor2_1 U58 ( .in0(v), .in1(n408), .out(net841));
inv1x_5 U59 ( .in0(e0), .out(net704));
inv1x_2 U60 ( .in0(net704), .out(net960));
nand3_4 U61 ( .in0(net702), .in1(net703), .in2(net704), .out(net970));
inv1x_2 U62 ( .in0(w), .out(net653));
nor2_2 U63 ( .in0(w), .in1(net685), .out(net689));
nor2_1 U64 ( .in0(w), .in1(net659), .out(net763));
inv1x_2 U65 ( .in0(net731), .out(net956));
inv1x_5 U66 ( .in0(c0), .out(net730));
nand3_4 U67 ( .in0(net732), .in1(net730), .in2(net894), .out(net897));
nand2_4 U68 ( .in0(net683), .in1(net730), .out(net729));
nand2_1 U69 ( .in0(net730), .in1(net674), .out(net758));
inv1x_13 U70 ( .in0(net701), .out(net1687));
nand4_3 U71 ( .in0(k), .in1(n512), .in2(n508), .in3(net674), .out(n410));
oai21_3 U72 ( .in0(i0), .in1(net699), .in2(net2956), .out(net896));
nand2_9 U73 ( .in0(v), .in1(net2959), .out(net936));
nand2_2 U74 ( .in0(net2959), .in1(net853), .out(net756));
nand2_4 U75 ( .in0(i0), .in1(net1620), .out(net2956));
inv1x_5 U76 ( .in0(net2959), .out(net776));
inv1x_2 U77 ( .in0(net680), .out(net2995));
inv1x_5 U78 ( .in0(net2994), .out(net924));
inv1x_4 U79 ( .in0(net2998), .out(net2857));
inv1x_8 U80 ( .in0(net680), .out(net2998));
aoi21_4 U81 ( .in0(net2956), .in1(net732), .in2(net1678), .out(net777));
aoi21_5 U82 ( .in0(net641), .in1(net642), .in2(net643), .out(n0));
oai22_2 U83 ( .in0(net742), .in1(n422), .in2(net742), .in3(n420), .out(net643));
inv1x_9 U84 ( .in0(n419), .out(n420));
aoi21_6 U85 ( .in0(net829), .in1(net830), .in2(n418), .out(n419));
oai21_3 U86 ( .in0(n416), .in1(net729), .in2(net827), .out(n418));
inv1x_13 U87 ( .in0(net687), .out(n416));
nor2_3 U88 ( .in0(n416), .in1(net758), .out(net759));
inv1x_2 U89 ( .in0(net739), .out(net829));
nand2_5 U90 ( .in0(n417), .in1(n421), .out(n422));
aoi22_1 U91 ( .in0(net830), .in1(net2857), .in2(n415), .in3(net830), .out(n421));
inv1x_2 U92 ( .in0(n413), .out(n415));
nand2_10 U93 ( .in0(n415), .in1(net741), .out(net739));
nand3_5 U94 ( .in0(n414), .in1(net738), .in2(d0), .out(n413));
inv1x_2 U95 ( .in0(v), .out(net691));
nand2_2 U96 ( .in0(net791), .in1(net691), .out(net843));
oai21_3 U97 ( .in0(n411), .in1(n412), .in2(v), .out(n414));
inv1x_3 U98 ( .in0(h0), .out(n412));
nor2_1 U99 ( .in0(o), .in1(z), .out(n411));
inv1x_3 U100 ( .in0(net686), .out(n417));
nor2_1 U101 ( .in0(d0), .in1(n417), .out(net813));
nor2_1 U102 ( .in0(net672), .in1(net673), .out(net671));
inv1x_3 U103 ( .in0(net867), .out(net672));
nor3_1 U104 ( .in0(net742), .in1(n423), .in2(n428), .out(net641));
nand3_4 U105 ( .in0(n429), .in1(net739), .in2(n430), .out(n428));
nand3_6 U106 ( .in0(n426), .in1(n432), .in2(n433), .out(n430));
nand3_3 U107 ( .in0(net936), .in1(net659), .in2(net924), .out(n433));
nand2_2 U108 ( .in0(j), .in1(n431), .out(n432));
nand2_2 U109 ( .in0(k), .in1(net648), .out(n431));
nor2_1 U110 ( .in0(net705), .in1(net703), .out(n426));
inv1x_9 U111 ( .in0(f0), .out(net703));
nand3_7 U112 ( .in0(net702), .in1(net703), .in2(net979), .out(net701));
inv1x_5 U113 ( .in0(h), .out(net705));
nand3_4 U114 ( .in0(net697), .in1(net705), .in2(net1592), .out(net865));
nand2_2 U115 ( .in0(n427), .in1(n425), .out(n429));
inv1x_5 U116 ( .in0(net682), .out(n425));
nand2_4 U117 ( .in0(net689), .in1(n425), .out(net688));
nor3_2 U118 ( .in0(net718), .in1(v), .in2(m), .out(n427));
inv1x_2 U119 ( .in0(c), .out(net718));
nand3_4 U120 ( .in0(net845), .in1(net944), .in2(net718), .out(net952));
aoi21_7 U121 ( .in0(net668), .in1(net669), .in2(n424), .out(n423));
nand3_5 U122 ( .in0(k0), .in1(net2857), .in2(net791), .out(n424));
nand2_2 U123 ( .in0(h), .in1(j0), .out(net795));
nand2_1 U124 ( .in0(h), .in1(f0), .out(net728));
nand2_10 U125 ( .in0(n434), .in1(net728), .out(net836));
nand2_4 U126 ( .in0(h), .in1(j0), .out(n434));
inv1x_3 U127 ( .in0(net774), .out(net1685));
inv1x_8 U128 ( .in0(net659), .out(net1681));
inv1x_8 U129 ( .in0(net1681), .out(net1682));
inv1x_2 U130 ( .in0(x), .out(net1678));
nand2_1 U131 ( .in0(n410), .in1(net709), .out(n435));
nor2_1 U132 ( .in0(net1592), .in1(net1668), .out(net788));
nand2_2 U133 ( .in0(net1620), .in1(net907), .out(net664));
nand2_9 U134 ( .in0(net1636), .in1(n436), .out(net894));
nand3_7 U135 ( .in0(net917), .in1(net1636), .in2(n436), .out(net741));
nand3_4 U136 ( .in0(i0), .in1(net1620), .in2(net679), .out(n436));
inv1x_3 U137 ( .in0(net1620), .out(net1668));
inv1x_9 U138 ( .in0(net1671), .out(net1592));
inv1x_5 U139 ( .in0(j0), .out(net1671));
nand3_5 U140 ( .in0(net830), .in1(net797), .in2(net3006), .out(net949));
nand3_3 U141 ( .in0(net748), .in1(net946), .in2(net904), .out(net669));
inv1x_8 U142 ( .in0(n435), .out(net904));
nand2_3 U143 ( .in0(n505), .in1(n504), .out(n437));
inv1x_2 U144 ( .in0(e0), .out(net979));
oai21_3 U145 ( .in0(net693), .in1(net688), .in2(net744), .out(n438));
nand2_2 U146 ( .in0(n491), .in1(n439), .out(n440));
inv1x_3 U147 ( .in0(n488), .out(n439));
inv1x_2 U148 ( .in0(n440), .out(n441));
inv1x_8 U149 ( .in0(net836), .out(net968));
inv1x_8 U150 ( .in0(net776), .out(net964));
inv1x_5 U151 ( .in0(net960), .out(net961));
aoi21_8 U152 ( .in0(n442), .in1(n443), .in2(c0), .out(p0));
aoi21_4 U153 ( .in0(k), .in1(net648), .in2(n445), .out(n444));
nor2_1 U154 ( .in0(v), .in1(u), .out(n446));
nor2_1 U155 ( .in0(net652), .in1(net653), .out(n447));
nor2_1 U156 ( .in0(b), .in1(net655), .out(n448));
aoi21_7 U157 ( .in0(n450), .in1(n451), .in2(net1682), .out(n449));
nor2_2 U158 ( .in0(net659), .in1(n453), .out(n452));
aoi21_4 U159 ( .in0(net664), .in1(net1636), .in2(n527), .out(n454));
inv1x_14 U160 ( .in0(n), .out(net674));
nand3_8 U161 ( .in0(n455), .in1(n456), .in2(net679), .out(net676));
nand3_2 U162 ( .in0(d0), .in1(net683), .in2(net684), .out(net682));
nand2_4 U163 ( .in0(net686), .in1(net687), .out(net685));
inv1x_5 U164 ( .in0(i0), .out(net697));
inv1x_2 U165 ( .in0(j0), .out(net699));
nand2_10 U166 ( .in0(h0), .in1(o), .out(net652));
inv1x_3 U167 ( .in0(k), .out(net707));
inv1x_2 U168 ( .in0(j), .out(net709));
inv1x_5 U169 ( .in0(g0), .out(net702));
inv1x_3 U170 ( .in0(m0), .out(n457));
nand2_11 U171 ( .in0(n458), .in1(n459), .out(net655));
nand2_1 U172 ( .in0(d0), .in1(net653), .out(net723));
inv1x_1 U173 ( .in0(x), .out(net679));
nand2_9 U174 ( .in0(net970), .in1(n460), .out(n453));
nand2_1 U175 ( .in0(z), .in1(h0), .out(net673));
inv1x_3 U176 ( .in0(b), .out(n461));
nand2_12 U177 ( .in0(n), .in1(o), .out(net686));
nand2_4 U178 ( .in0(n463), .in1(net748), .out(n462));
nand2_2 U179 ( .in0(n464), .in1(net709), .out(net749));
oai22_3 U180 ( .in0(n446), .in1(net723), .in2(net754), .in3(n453), .out(n465));
nor2_2 U181 ( .in0(d0), .in1(net652), .out(n466));
nand2_2 U182 ( .in0(j), .in1(net699), .out(n445));
nor2_4 U183 ( .in0(c), .in1(f), .out(n459));
nor2_5 U184 ( .in0(e), .in1(g), .out(n458));
nor2_1 U185 ( .in0(n448), .in1(net961), .out(n467));
nor2_1 U186 ( .in0(net765), .in1(net766), .out(n468));
oai21_3 U187 ( .in0(n444), .in1(net968), .in2(n468), .out(n469));
aoi21_7 U188 ( .in0(n467), .in1(n471), .in2(n457), .out(n470));
aoi21_7 U189 ( .in0(n473), .in1(n474), .in2(n469), .out(n472));
nand2_2 U190 ( .in0(net686), .in1(net687), .out(n475));
aoi21_4 U191 ( .in0(x), .in1(net970), .in2(net774), .out(n450));
nor2_2 U192 ( .in0(net754), .in1(net776), .out(n476));
nor2_2 U193 ( .in0(net783), .in1(n438), .out(n442));
aoi21_9 U194 ( .in0(n472), .in1(n470), .in2(n477), .out(n443));
aoi21_1 U195 ( .in0(net777), .in1(n476), .in2(n452), .out(n478));
nand3_4 U196 ( .in0(n479), .in1(n480), .in2(n478), .out(n477));
nand3_3 U197 ( .in0(net961), .in1(net2857), .in2(net652), .out(n481));
nand2_2 U198 ( .in0(l0), .in1(net791), .out(n482));
nor2_2 U199 ( .in0(n481), .in1(n482), .out(n483));
nor2_1 U200 ( .in0(net729), .in1(net685), .out(net799));
nor2_2 U201 ( .in0(net707), .in1(n461), .out(n484));
aoi21_4 U202 ( .in0(b), .in1(j), .in2(r), .out(n485));
nor2_1 U203 ( .in0(a), .in1(u), .out(n486));
nor2_1 U204 ( .in0(f), .in1(e), .out(n487));
nand2_2 U205 ( .in0(n487), .in1(n486), .out(n488));
nand2_2 U206 ( .in0(net686), .in1(n490), .out(n489));
nor2_2 U207 ( .in0(n489), .in1(net682), .out(n491));
nor2_1 U208 ( .in0(net729), .in1(net655), .out(n492));
nand2_2 U209 ( .in0(net791), .in1(net1685), .out(n493));
nor2_1 U210 ( .in0(n495), .in1(n493), .out(n494));
nand2_2 U211 ( .in0(l0), .in1(n434), .out(n495));
aoi21_10 U212 ( .in0(n496), .in1(n494), .in2(net824), .out(net645));
nor2_2 U213 ( .in0(net836), .in1(n497), .out(n463));
aoi21_4 U214 ( .in0(n498), .in1(n499), .in2(n454), .out(net668));
nor2_2 U215 ( .in0(j), .in1(net655), .out(n500));
nand2_2 U216 ( .in0(k0), .in1(n434), .out(n501));
nor2_1 U217 ( .in0(n501), .in1(net843), .out(net845));
nor2_2 U218 ( .in0(v), .in1(net2857), .out(n502));
aoi21_7 U219 ( .in0(net841), .in1(d0), .in2(net774), .out(n503));
inv1x_6 U220 ( .in0(l), .out(n504));
inv1x_3 U221 ( .in0(t), .out(n505));
inv1x_6 U222 ( .in0(s), .out(n506));
inv1x_15 U223 ( .in0(b0), .out(n455));
inv1x_15 U224 ( .in0(q), .out(n456));
inv1x_3 U225 ( .in0(g), .out(n490));
nand2_2 U226 ( .in0(net853), .in1(net867), .out(net866));
nand3_9 U227 ( .in0(net956), .in1(net2857), .in2(n507), .out(net827));
inv1x_3 U228 ( .in0(n462), .out(n498));
nand2_11 U229 ( .in0(m), .in1(r), .out(net687));
inv1x_2 U230 ( .in0(net701), .out(net732));
nand4_4 U231 ( .in0(n456), .in1(n455), .in2(net687), .in3(net686), .out(n460));
nand2_2 U232 ( .in0(n505), .in1(n504), .out(n508));
nand3_4 U233 ( .in0(n437), .in1(net674), .in2(n517), .out(net648));
inv1x_2 U234 ( .in0(net652), .out(net774));
inv1x_9 U235 ( .in0(net676), .out(net683));
oai21_3 U236 ( .in0(net676), .in1(n475), .in2(net754), .out(n451));
inv1x_6 U237 ( .in0(net655), .out(net748));
nand2_11 U238 ( .in0(i), .in1(g0), .out(net791));
inv1x_3 U239 ( .in0(net791), .out(net766));
inv1x_3 U240 ( .in0(net673), .out(net765));
nand3_4 U241 ( .in0(net683), .in1(net896), .in2(net759), .out(n509));
nand2_10 U242 ( .in0(net897), .in1(n509), .out(n510));
nand2_6 U243 ( .in0(n466), .in1(n510), .out(net744));
nand2_2 U244 ( .in0(b), .in1(m), .out(n511));
inv1x_3 U245 ( .in0(n511), .out(n497));
nand4_5 U246 ( .in0(k), .in1(n512), .in2(n508), .in3(net674), .out(n464));
nand2_2 U247 ( .in0(m), .in1(n435), .out(n513));
nand2_2 U248 ( .in0(net748), .in1(n513), .out(n471));
nand2_9 U249 ( .in0(net664), .in1(net865), .out(n499));
nand2_2 U250 ( .in0(m), .in1(net749), .out(n514));
nand2_2 U251 ( .in0(c), .in1(n514), .out(n515));
nand2_2 U252 ( .in0(net763), .in1(n515), .out(n474));
inv1x_3 U253 ( .in0(n449), .out(n480));
oai21_2 U254 ( .in0(n447), .in1(n465), .in2(net964), .out(n479));
nand2_2 U255 ( .in0(v), .in1(d0), .out(net911));
nand4_3 U256 ( .in0(n437), .in1(net674), .in2(n484), .in3(n517), .out(n516));
nand2_1 U257 ( .in0(n485), .in1(n516), .out(n518));
nand2_1 U258 ( .in0(m), .in1(n518), .out(n519));
nand2_2 U259 ( .in0(net986), .in1(net1678), .out(n520));
nand3_6 U260 ( .in0(net917), .in1(net865), .in2(n520), .out(n507));
nand2_9 U261 ( .in0(net788), .in1(net907), .out(n521));
nand2_1 U262 ( .in0(net920), .in1(n521), .out(n522));
nand2_2 U263 ( .in0(n441), .in1(n519), .out(n523));
nand4_3 U264 ( .in0(n492), .in1(n522), .in2(net813), .in3(n519), .out(n524));
nand3_4 U265 ( .in0(n523), .in1(net827), .in2(n524), .out(n496));
nand2_4 U266 ( .in0(net1682), .in1(net924), .out(net867));
nand2_1 U267 ( .in0(n483), .in1(n522), .out(net927));
nand2_1 U268 ( .in0(net765), .in1(net867), .out(net928));
nand3_2 U269 ( .in0(net830), .in1(net825), .in2(net741), .out(net743));
nand2_1 U270 ( .in0(n500), .in1(n526), .out(n525));
nand2_10 U271 ( .in0(net968), .in1(net961), .out(n527));
nand3_4 U272 ( .in0(n527), .in1(n462), .in2(n525), .out(net944));
nand3_5 U273 ( .in0(n521), .in1(net865), .in2(net945), .out(net946));
inv1x_2 U274 ( .in0(net728), .out(net853));
nand2_2 U275 ( .in0(n499), .in1(net2857), .out(n473));
nand2_9 U276 ( .in0(d), .in1(n506), .out(n517));
inv1x_3 U277 ( .in0(net949), .out(net824));
nand2_4 U278 ( .in0(d), .in1(n506), .out(n512));
nand4_5 U279 ( .in0(k), .in1(n512), .in2(n437), .in3(net674), .out(n526));
nand3_4 U280 ( .in0(n528), .in1(net952), .in2(n503), .out(net852));
nand3_5 U281 ( .in0(n502), .in1(net904), .in2(c), .out(n528));
endmodule
