VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

LAYER nwell
  TYPE  MASTERSLICE ;
END nwell

LAYER nselect
  TYPE  MASTERSLICE ;
END nselect

LAYER pselect
  TYPE  MASTERSLICE ;
END pselect

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cp
  TYPE	CUT ;
  SPACING	0.3 ;
END cp

LAYER ca
  TYPE	CUT ;
  SPACING	0.3 ;
END ca

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.8  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0 ;
  CAPACITANCE	CPERSQDIST 0 ;
  CURRENTDEN 0 ;
END metal1

LAYER via
  TYPE	CUT ;
  SPACING	0.3 ;
END via

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.8  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0 ;
  CAPACITANCE	CPERSQDIST 0 ;
  CURRENTDEN 0 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.3 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.8  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  RESISTANCE	RPERSQ 0 ;
  CAPACITANCE	CPERSQDIST 0 ;
  CURRENTDEN 0 ;
END metal3

LAYER LAYER42
  TYPE	MASTERSLICE ;
END LAYER42

LAYER LAYER44
  TYPE	MASTERSLICE ;
END LAYER44

LAYER LAYER45
  TYPE	MASTERSLICE ;
END LAYER45

LAYER text
  TYPE	VIRTUAL ;
END text

SPACING
  SAMENET metal1  metal1	0.3 ;
  SAMENET metal2  metal2	0.3 ;
  SAMENET metal3  metal3	0.3 ;
  SAMENET ca  ca	0.3 ;
  SAMENET ca  cp	0.3 ;
  SAMENET cp  cp	0.3 ;
  SAMENET ca  via	0.3 ;
  SAMENET cp  via	0.3 ;
  SAMENET via  via	0.3 ;
  SAMENET via2  via2	0.3 ;
  SAMENET via  via2	0.3 ;
END SPACING

VIA PTAP DEFAULT
  LAYER pactive ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER ca ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END PTAP

VIA NTAP DEFAULT
  LAYER nactive ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER ca ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END NTAP

VIA M1_POLY DEFAULT
  LAYER poly ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER cp ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M1_POLY

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER via ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER via2 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END M3_M2


VIARULE VIAGEN12 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via ;
    RECT -0.10 -0.10 0.10 0.10 ;
    SPACING 0.8 BY 0.8 ;
END VIAGEN12

VIARULE VIAGEN23 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.10 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
    RECT -0.10 -0.10 0.10 0.10 ;
    SPACING 0.8 BY 0.8 ;
END VIAGEN23

VIARULE Turn1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END Turn1

VIARULE Turn2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END Turn2

VIARULE Turn3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END Turn3

SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SIZE        8.000 BY 118.000 ;
END  CoreSite

SITE  TDCoverSite
    CLASS       CORE ;
    SIZE        1.000 BY 1.000 ;
END  TDCoverSite

SITE  SBlockSite
    CLASS       CORE ;
    SIZE        1.000 BY 1.000 ;
END  SBlockSite

SITE  PortCellSite
    CLASS       PAD ;
    SIZE        1.000 BY 1.000 ;
END  PortCellSite

SITE  Core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SIZE        8.000 BY 118.000 ;
END  Core

MACRO invload
  CLASS CORE ;
  FOREIGN invload -0.360 -2.270 ;
  ORIGIN 0.360 2.270 ;
  SIZE 11.520 BY 5.040 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -0.360 2.370 11.160 3.170 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -0.360 -2.670 11.160 -1.870 ;
    END
  END gnd!
  PIN out
    DIRECTION OUTPUT ;
    PORT
    LAYER METAL2 ;
    RECT 0.580 -0.140 0.865 0.240 ;
    END
  END out
  PIN in0
    DIRECTION INPUT ;
    PORT
    LAYER METAL2 ;
    RECT -0.140 -0.140 0.140 0.240 ;
    END
  END in0
  OBS
    LAYER NWELL ;
    RECT -0.790 0.000 11.590 3.310 ;
    LAYER NINP ;
    RECT -0.390 -1.725 11.190 0.000 ;
    RECT -0.460 2.225 11.260 2.990 ;
    LAYER PINP ;
    RECT -0.390 0.000 11.190 2.225 ;
    RECT -0.460 -2.490 11.260 -1.725 ;
    LAYER N2V ;
    RECT -0.390 -1.725 11.190 0.000 ;
    LAYER P2V ;
    RECT -0.390 0.000 11.190 2.225 ;
    LAYER DIFF ;
    RECT -0.360 2.325 11.160 2.880 ;
    RECT -0.210 -1.370 11.010 -0.435 ;
    RECT -0.360 -2.380 11.160 -1.825 ;
    RECT -0.210 0.450 11.010 1.855 ;
    LAYER POLY1 ;
    RECT 0.270 0.000 0.450 2.075 ;
    RECT 0.990 0.000 1.170 2.075 ;
    RECT 0.270 -0.330 0.990 0.330 ;
    RECT 1.710 0.000 1.890 2.075 ;
    RECT 0.990 -0.330 1.710 0.330 ;
    RECT 2.430 0.000 2.610 2.075 ;
    RECT 1.710 -0.330 2.430 0.330 ;
    RECT 3.150 0.000 3.330 2.075 ;
    RECT 2.430 -0.330 3.150 0.330 ;
    RECT 3.870 0.000 4.050 2.075 ;
    RECT 3.150 -0.330 3.870 0.330 ;
    RECT 4.590 0.000 4.770 2.075 ;
    RECT 3.870 -0.330 4.590 0.330 ;
    RECT 5.310 0.000 5.490 2.075 ;
    RECT 4.590 -0.330 5.310 0.330 ;
    RECT 6.030 0.000 6.210 2.075 ;
    RECT 5.310 -0.330 6.030 0.330 ;
    RECT 6.750 0.000 6.930 2.075 ;
    RECT 6.030 -0.330 6.750 0.330 ;
    RECT 7.470 0.000 7.650 2.075 ;
    RECT 6.750 -0.330 7.470 0.330 ;
    RECT 8.190 0.000 8.370 2.075 ;
    RECT 7.470 -0.330 8.190 0.330 ;
    RECT 8.910 0.000 9.090 2.075 ;
    RECT 8.190 -0.330 8.910 0.330 ;
    RECT 9.630 0.000 9.810 2.075 ;
    RECT 8.910 -0.330 9.630 0.330 ;
    RECT 10.350 0.000 10.530 2.075 ;
    RECT 9.630 -0.330 10.350 0.330 ;
    RECT 0.270 -1.590 0.450 0.000 ;
    RECT 0.990 -1.590 1.170 0.000 ;
    RECT 0.270 -0.330 0.990 0.330 ;
    RECT 1.710 -1.590 1.890 0.000 ;
    RECT 0.990 -0.330 1.710 0.330 ;
    RECT 2.430 -1.590 2.610 0.000 ;
    RECT 1.710 -0.330 2.430 0.330 ;
    RECT 3.150 -1.590 3.330 0.000 ;
    RECT 2.430 -0.330 3.150 0.330 ;
    RECT 3.870 -1.590 4.050 0.000 ;
    RECT 3.150 -0.330 3.870 0.330 ;
    RECT 4.590 -1.590 4.770 0.000 ;
    RECT 3.870 -0.330 4.590 0.330 ;
    RECT 5.310 -1.590 5.490 0.000 ;
    RECT 4.590 -0.330 5.310 0.330 ;
    RECT 6.030 -1.590 6.210 0.000 ;
    RECT 5.310 -0.330 6.030 0.330 ;
    RECT 6.750 -1.590 6.930 0.000 ;
    RECT 6.030 -0.330 6.750 0.330 ;
    RECT 7.470 -1.590 7.650 0.000 ;
    RECT 6.750 -0.330 7.470 0.330 ;
    RECT 8.190 -1.590 8.370 0.000 ;
    RECT 7.470 -0.330 8.190 0.330 ;
    RECT 8.910 -1.590 9.090 0.000 ;
    RECT 8.190 -0.330 8.910 0.330 ;
    RECT 9.630 -1.590 9.810 0.000 ;
    RECT 8.910 -0.330 9.630 0.330 ;
    RECT 10.350 -1.590 10.530 0.000 ;
    RECT 9.630 -0.330 10.350 0.330 ;
    RECT -0.020 -0.130 0.400 0.290 ;
    LAYER METAL1 ;
    RECT -0.360 2.370 11.160 3.170 ;
    RECT -0.360 -2.670 11.160 -1.870 ;
    RECT -0.190 -0.090 0.305 0.325 ;
    RECT 0.535 -0.090 0.915 0.190 ;
    RECT -0.170 1.035 0.170 1.265 ;
    RECT -0.115 1.150 0.115 2.770 ;
    RECT 0.550 1.035 0.890 1.265 ;
    RECT 0.605 0.000 0.835 1.150 ;
    RECT 1.270 1.035 1.610 1.265 ;
    RECT 1.325 1.150 1.555 2.770 ;
    RECT 1.990 1.035 2.330 1.265 ;
    RECT 2.045 0.000 2.275 1.150 ;
    RECT 0.720 -0.090 2.160 0.140 ;
    RECT 2.710 1.035 3.050 1.265 ;
    RECT 2.765 1.150 2.995 2.770 ;
    RECT 3.430 1.035 3.770 1.265 ;
    RECT 3.485 0.000 3.715 1.150 ;
    RECT 2.160 -0.090 3.600 0.140 ;
    RECT 4.150 1.035 4.490 1.265 ;
    RECT 4.205 1.150 4.435 2.770 ;
    RECT 4.870 1.035 5.210 1.265 ;
    RECT 4.925 0.000 5.155 1.150 ;
    RECT 3.600 -0.090 5.040 0.140 ;
    RECT 5.590 1.035 5.930 1.265 ;
    RECT 5.645 1.150 5.875 2.770 ;
    RECT 6.310 1.035 6.650 1.265 ;
    RECT 6.365 0.000 6.595 1.150 ;
    RECT 5.040 -0.090 6.480 0.140 ;
    RECT 7.030 1.035 7.370 1.265 ;
    RECT 7.085 1.150 7.315 2.770 ;
    RECT 7.750 1.035 8.090 1.265 ;
    RECT 7.805 0.000 8.035 1.150 ;
    RECT 6.480 -0.090 7.920 0.140 ;
    RECT 8.470 1.035 8.810 1.265 ;
    RECT 8.525 1.150 8.755 2.770 ;
    RECT 9.190 1.035 9.530 1.265 ;
    RECT 9.245 0.000 9.475 1.150 ;
    RECT 7.920 -0.090 9.360 0.140 ;
    RECT 9.910 1.035 10.250 1.265 ;
    RECT 9.965 1.150 10.195 2.770 ;
    RECT 10.630 1.035 10.970 1.265 ;
    RECT 10.685 0.000 10.915 1.150 ;
    RECT 9.360 -0.090 10.800 0.140 ;
    RECT -0.170 -1.020 0.170 -0.790 ;
    RECT -0.115 -2.270 0.115 -0.905 ;
    RECT 0.550 -1.020 0.890 -0.790 ;
    RECT 0.605 -0.905 0.835 0.000 ;
    RECT 1.270 -1.020 1.610 -0.790 ;
    RECT 1.325 -2.270 1.555 -0.905 ;
    RECT 1.990 -1.020 2.330 -0.790 ;
    RECT 2.045 -0.905 2.275 0.000 ;
    RECT 0.720 -0.090 2.160 0.140 ;
    RECT 2.710 -1.020 3.050 -0.790 ;
    RECT 2.765 -2.270 2.995 -0.905 ;
    RECT 3.430 -1.020 3.770 -0.790 ;
    RECT 3.485 -0.905 3.715 0.000 ;
    RECT 2.160 -0.090 3.600 0.140 ;
    RECT 4.150 -1.020 4.490 -0.790 ;
    RECT 4.205 -2.270 4.435 -0.905 ;
    RECT 4.870 -1.020 5.210 -0.790 ;
    RECT 4.925 -0.905 5.155 0.000 ;
    RECT 3.600 -0.090 5.040 0.140 ;
    RECT 5.590 -1.020 5.930 -0.790 ;
    RECT 5.645 -2.270 5.875 -0.905 ;
    RECT 6.310 -1.020 6.650 -0.790 ;
    RECT 6.365 -0.905 6.595 0.000 ;
    RECT 5.040 -0.090 6.480 0.140 ;
    RECT 7.030 -1.020 7.370 -0.790 ;
    RECT 7.085 -2.270 7.315 -0.905 ;
    RECT 7.750 -1.020 8.090 -0.790 ;
    RECT 7.805 -0.905 8.035 0.000 ;
    RECT 6.480 -0.090 7.920 0.140 ;
    RECT 8.470 -1.020 8.810 -0.790 ;
    RECT 8.525 -2.270 8.755 -0.905 ;
    RECT 9.190 -1.020 9.530 -0.790 ;
    RECT 9.245 -0.905 9.475 0.000 ;
    RECT 7.920 -0.090 9.360 0.140 ;
    RECT 9.910 -1.020 10.250 -0.790 ;
    RECT 9.965 -2.270 10.195 -0.905 ;
    RECT 10.630 -1.020 10.970 -0.790 ;
    RECT 10.685 -0.905 10.915 0.000 ;
    RECT 9.360 -0.090 10.800 0.140 ;
    LAYER CONT ;
    RECT 0.080 -0.030 0.300 0.190 ;
    RECT -0.110 2.425 0.110 2.645 ;
    RECT -0.110 -2.145 0.110 -1.925 ;
    RECT 0.610 2.425 0.830 2.645 ;
    RECT 0.610 -2.145 0.830 -1.925 ;
    RECT 1.330 2.425 1.550 2.645 ;
    RECT 1.330 -2.145 1.550 -1.925 ;
    RECT 2.050 2.425 2.270 2.645 ;
    RECT 2.050 -2.145 2.270 -1.925 ;
    RECT 2.770 2.425 2.990 2.645 ;
    RECT 2.770 -2.145 2.990 -1.925 ;
    RECT 3.490 2.425 3.710 2.645 ;
    RECT 3.490 -2.145 3.710 -1.925 ;
    RECT 4.210 2.425 4.430 2.645 ;
    RECT 4.210 -2.145 4.430 -1.925 ;
    RECT 4.930 2.425 5.150 2.645 ;
    RECT 4.930 -2.145 5.150 -1.925 ;
    RECT 5.650 2.425 5.870 2.645 ;
    RECT 5.650 -2.145 5.870 -1.925 ;
    RECT 6.370 2.425 6.590 2.645 ;
    RECT 6.370 -2.145 6.590 -1.925 ;
    RECT 7.090 2.425 7.310 2.645 ;
    RECT 7.090 -2.145 7.310 -1.925 ;
    RECT 7.810 2.425 8.030 2.645 ;
    RECT 7.810 -2.145 8.030 -1.925 ;
    RECT 8.530 2.425 8.750 2.645 ;
    RECT 8.530 -2.145 8.750 -1.925 ;
    RECT 9.250 2.425 9.470 2.645 ;
    RECT 9.250 -2.145 9.470 -1.925 ;
    RECT 9.970 2.425 10.190 2.645 ;
    RECT 9.970 -2.145 10.190 -1.925 ;
    RECT 10.690 2.425 10.910 2.645 ;
    RECT 10.690 -2.145 10.910 -1.925 ;
    RECT -0.110 1.040 0.110 1.260 ;
    RECT 0.610 1.040 0.830 1.260 ;
    RECT 1.330 1.040 1.550 1.260 ;
    RECT 2.050 1.040 2.270 1.260 ;
    RECT 2.770 1.040 2.990 1.260 ;
    RECT 3.490 1.040 3.710 1.260 ;
    RECT 4.210 1.040 4.430 1.260 ;
    RECT 4.930 1.040 5.150 1.260 ;
    RECT 5.650 1.040 5.870 1.260 ;
    RECT 6.370 1.040 6.590 1.260 ;
    RECT 7.090 1.040 7.310 1.260 ;
    RECT 7.810 1.040 8.030 1.260 ;
    RECT 8.530 1.040 8.750 1.260 ;
    RECT 9.250 1.040 9.470 1.260 ;
    RECT 9.970 1.040 10.190 1.260 ;
    RECT 10.690 1.040 10.910 1.260 ;
    RECT -0.110 -1.015 0.110 -0.785 ;
    RECT 0.610 -1.015 0.830 -0.785 ;
    RECT 1.330 -1.015 1.550 -0.785 ;
    RECT 2.050 -1.015 2.270 -0.785 ;
    RECT 2.770 -1.015 2.990 -0.785 ;
    RECT 3.490 -1.015 3.710 -0.785 ;
    RECT 4.210 -1.015 4.430 -0.785 ;
    RECT 4.930 -1.015 5.150 -0.785 ;
    RECT 5.650 -1.015 5.870 -0.785 ;
    RECT 6.370 -1.015 6.590 -0.785 ;
    RECT 7.090 -1.015 7.310 -0.785 ;
    RECT 7.810 -1.015 8.030 -0.785 ;
    RECT 8.530 -1.015 8.750 -0.785 ;
    RECT 9.250 -1.015 9.470 -0.785 ;
    RECT 9.970 -1.015 10.190 -0.785 ;
    RECT 10.690 -1.015 10.910 -0.785 ;
    LAYER VIA12 ;
    RECT -0.130 -0.080 0.130 0.180 ;
    RECT 0.595 -0.080 0.855 0.180 ;
  END
END invload
MACRO filler
  CLASS CORE ;
  FOREIGN filler -20.000 -56.000 ;
  ORIGIN 20.000 56.000 ;
  SIZE 16.000 BY 112.000 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -20.000 54.000 -4.000 58.000 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
    LAYER METAL1 ;
    RECT -20.000 -58.000 -4.000 -54.000 ;
    END
  END gnd!
  PIN shield_0
    DIRECTION INOUT ;
    PORT
    LAYER METAL2 ;
    RECT -6.000 -58.000 -2.000 58.000 ;
    END
  END shield_0
  PIN shield_1
    DIRECTION INOUT ;
    PORT
    LAYER METAL2 ;
    RECT -22.000 -58.000 -18.000 58.000 ;
    END
  END shield_1
  OBS
    LAYER NWELL ;
    RECT -24.000 0.000 0.000 62.000 ;
    LAYER NIMP ;
    RECT -20.000 52.000 -4.000 60.000 ;
    RECT -20.000 -52.000 -4.000 0.000 ;
    LAYER PIMP ;
    RECT -20.000 -60.000 -4.000 -52.000 ;
    RECT -20.000 0.000 -4.000 52.000 ;
    LAYER DIFF ;
    RECT -18.000 54.000 -6.000 58.000 ;
    LAYER DIFF ;
    RECT -18.000 -58.000 -6.000 -54.000 ;
    LAYER CONT ;
    RECT -9.000 55.000 -7.000 57.000 ;
    RECT -9.000 -57.000 -7.000 -55.000 ;
    RECT -17.000 55.000 -15.000 57.000 ;
    RECT -17.000 -57.000 -15.000 -55.000 ;
  END
END filler
END LIBRARY
